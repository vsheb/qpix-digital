    .INIT_00(256'h022ffd250002f013022ffd2072a0b002022ffd2072a2f01f022ffd2072a01004),
    .INIT_01(256'h022ffd20700206dc022ffd3680b32208022ffd1d0001d002022ffd0b0320b032),
    .INIT_02(256'h022ffd25000324f1022ffd206dc1d001022ffd2071e0b032022ffd207182078c),
    .INIT_03(256'h022ffd206dc2074d022ffd206fc01004022ffd20712324f1022ffd207001d002),
    .INIT_04(256'h022ffd368182f03a022ffd1d00011001022ffd0b0320b03a022ffd2500022008),
    .INIT_05(256'h022ffd206dc1f000022ffd207020b017022ffd207161d000022ffd207040b016),
    .INIT_06(256'h022ffd207001f000022ffd207000b019022ffd207041f000022ffd250000b018),
    .INIT_07(256'h022ffd206fc1f000022ffd2071a0b01b022ffd207e91f000022ffd206dc0b01a),
    .INIT_08(256'h022ffd0b00f1f000022ffd141060b01d022ffd0b1131f000022ffd206de0b01c),
    .INIT_09(256'h022ffd206bd1d001022ffd206bd0b032022ffd00c00208a5022ffd0401036017),
    .INIT_0A(256'h022ffd206b522008022ffd0b00e324cd022ffd207301d002022ffd206c73247a),
    .INIT_0B(256'h022ffd206b50be11022ffd0b00c0bd10022ffd206b52f01e022ffd0b00d01001),
    .INIT_0C(256'h022ffd206de13f00022ffd206fc13e00022ffd2071211d01022ffd206dc0bf12),
    .INIT_0D(256'h022ffd0b0122ff12022ffd1410603f01022ffd0b1132fe11022ffd206e82fd10),
    .INIT_0E(256'h022ffd206b52f00f022ffd0b01103001022ffd206b50b00f022ffd0401020b5f),
    .INIT_0F(256'h022ffd2500003e7e022ffd206dc0be0e022ffd206b50307e022ffd0b0100b03b),
    .INIT_10(256'h022ffd0bc1620911022ffd3487e208fa022ffd1dcff3625d022ffd0bc171c0e0),
    .INIT_11(256'h022ffd1dcff1f000022ffd0bc190b017022ffd348841d000022ffd1dcff0b016),
    .INIT_12(256'h022ffd348841f000022ffd1dcff0b019022ffd0bc181f000022ffd3487e0b018),
    .INIT_13(256'h022ffd0bc1a1f000022ffd3487e0b01b022ffd1dcff1f000022ffd0bc1b0b01a),
    .INIT_14(256'h022ffd1dcff1f000022ffd0bc1d0b01d022ffd348841f000022ffd1dcff0b01c),
    .INIT_15(256'h022ffd348842077b022ffd1dcff2075c022ffd0bc1c2225d022ffd3487e36256),
    .INIT_16(256'h022ffd328622074d022ffd1dd0001004022ffd0bd202078c022ffd25000206dc),
    .INIT_17(256'h022ffd2088a2b40f022ffd0bc162b20f022ffd2087e208a5022ffd0bc1722008),
    .INIT_18(256'h022ffd1dd002077b022ffd0bd212074d022ffd2089001002022ffd0bc202b80f),
    .INIT_19(256'h022ffd0bc180900e022ffd2087e2f032022ffd0bc1901000022ffd3286b22008),
    .INIT_1A(256'h022ffd0bd222f007022ffd2089009017022ffd0bc2132296022ffd2088a0d004),
    .INIT_1B(256'h022ffd2087e2f009022ffd0bc1b09019022ffd328742f008022ffd1dd0009018),
    .INIT_1C(256'h022ffd208902f00b022ffd0bc220901b022ffd2088a2f00a022ffd0bc1a0901a),
    .INIT_1D(256'h022ffd0bc1d3627c022ffd3287d1d0a0022ffd1dd00030f0022ffd0bd232b04e),
    .INIT_1E(256'h022ffd0bc23223ef022ffd2088a323ee022ffd0bc1c0d002022ffd2087e09002),
    .INIT_1F(256'h022ffd207021d0b0022ffd20728223ee022ffd250003627f022ffd208901d0e0),
    .INIT_20(256'h022ffd250002dc01022ffd206de03c0f022ffd206b60bc07022ffd206de36289),
    .INIT_21(256'h022ffd206b6206dc022ffd206de206b6022ffd20722206de022ffd206fe2071e),
    .INIT_22(256'h022ffd2072220724022ffd206fe3628d022ffd250001d0d0022ffd206dc22003),
    .INIT_23(256'h022ffd2500020702022ffd206de36291022ffd206b61d0f0022ffd206de2240b),
    .INIT_24(256'h022ffd206b60d080022ffd206de32414022ffd207261d0c0022ffd20712223fb),
    .INIT_25(256'h022ffd2b00a0d020022ffd2b0090900d022ffd25000223ec022ffd206dc32414),
    .INIT_26(256'h022ffd01c00362a0022ffd209091d04f022ffd2b08e09006022ffd2b1bb363ee),
    .INIT_27(256'h022ffd01c10223ef022ffd25000323ee022ffd200590d002022ffd208ae09002),
    .INIT_28(256'h022ffd208ae206dc022ffd01c0720720022ffd25000362a7022ffd208ae1d053),
    .INIT_29(256'h022ffd250001d052022ffd208ae223ed022ffd01c0d20793022ffd2500020784),
    .INIT_2A(256'h022ffd01c0409006022ffd2500020733022ffd208ae2071e022ffd01c01362be),
    .INIT_2B(256'h022ffd01e0020733022ffd01d00206de022ffd25000363ec022ffd208ae1d020),
    .INIT_2C(256'h022ffd01100206e8022ffd01080363ec022ffd208dd1d030022ffd01f0009006),
    .INIT_2D(256'h022ffd2b3893a3ec022ffd25000206a9022ffd208bd09006022ffd208d420733),
    .INIT_2E(256'h022ffd2090920730022ffd2b08e206c7022ffd2b63b00100022ffd2b00a2d001),
    .INIT_2F(256'h022ffd2b37b362c2022ffd2b00a1d055022ffd2b1c922003022ffd25000206dc),
    .INIT_30(256'h022ffd2b649362c6022ffd250001d044022ffd209092240b022ffd2b08e20724),
    .INIT_31(256'h022ffd20909362d7022ffd2b08e1d04e022ffd2b0bb223fb022ffd2b72a20702),
    .INIT_32(256'h022ffd2b57b1d020022ffd2b20a09006022ffd2b64920733022ffd2500020716),
    .INIT_33(256'h022ffd2b20a206cc022ffd2b6c90120a022ffd20909206de022ffd2b08e363ec),
    .INIT_34(256'h022ffd250002fc09022ffd209092fb08022ffd2b08e2fa07022ffd2b63b3a3ec),
    .INIT_35(256'h022ffd2d1081d054022ffd2d00822420022ffd2b4192fe0b022ffd2b00a2fd0a),
    .INIT_36(256'h022ffd2d10809006022ffd2d00820733022ffd2b25920722022ffd2b00a3632a),
    .INIT_37(256'h022ffd2dc080120a022ffd2b289206de022ffd2b00a363ec022ffd250001d020),
    .INIT_38(256'h022ffd250002fb3f022ffd2df082fa3e022ffd2de083a3ec022ffd2dd08206cc),
    .INIT_39(256'h022ffd09d08322e9022ffd09c080de80022ffd2b28932308022ffd2b00a1dec0),
    .INIT_3A(256'h022ffd208b7206a2022ffd25000206a2022ffd09f08206a2022ffd09e08223ec),
    .INIT_3B(256'h022ffd208bd206a2022ffd208dd363ec022ffd2500018fa0022ffd208e40ba02),
    .INIT_3C(256'h022ffd208d42ff0f022ffd011002fe0e022ffd010202fd0d022ffd250002fc0c),
    .INIT_3D(256'h022ffd0bc0c0be11022ffd0bd0d0bd10022ffd0be0e206dc022ffd0bf0f20aad),
    .INIT_3E(256'h022ffd208ab206b6022ffd208f100cf0022ffd2500020700022ffd208ee0bf12),
    .INIT_3F(256'h022ffd25000206b6022ffd2090000cd0022ffd25000206b6022ffd208c300ce0),
    .INIT_40(256'h022ffd208d4206c7022ffd01101206bd022ffd01080206bd022ffd208f10bc3f),
    .INIT_41(256'h022ffd208c9223ec022ffd208a8206b6022ffd208bd0bc3e022ffd208b720730),
    .INIT_42(256'h022ffd369090ba02022ffd0d008206a2022ffd0900e206a2022ffd25000206a2),
    .INIT_43(256'h022ffd3290d2fc10022ffd0d002206a2022ffd0900e363ec022ffd2500018ea0),
    .INIT_44(256'h022ffd2f116206dc022ffd0110020b5f022ffd370012fe12022ffd250002fd11),
    .INIT_45(256'h022ffd2f11a0bc0f022ffd2f1190bd0e022ffd2f1180be0d022ffd2f1170bf0c),
    .INIT_46(256'h022ffd0108420730022ffd2f11d206c7022ffd2f11c206bd022ffd2f11b206bd),
    .INIT_47(256'h022ffd11001206b6022ffd2b00b00ce0022ffd2b00a206b6022ffd2b6c900cd0),
    .INIT_48(256'h022ffd1d0ff206bd022ffd209860bc3f022ffd2092c206b6022ffd2092700cf0),
    .INIT_49(256'h022ffd09c080bc3e022ffd2500020730022ffd37000206c7022ffd3691f206bd),
    .INIT_4A(256'h022ffd2500036348022ffd09f081d058022ffd09e08223ec022ffd09d08206b6),
    .INIT_4B(256'h022ffd329572072a022ffd1d0c23e348022ffd329420d004022ffd1d0c109002),
    .INIT_4C(256'h022ffd20975363ec022ffd001e01d020022ffd2097509006022ffd001f020733),
    .INIT_4D(256'h022ffd209753a3ec022ffd001c0206cc022ffd2097501208022ffd001d0206de),
    .INIT_4E(256'h022ffd2f12c2fc36022ffd2f12a2fb35022ffd2f1282fa34022ffd01100206dc),
    .INIT_4F(256'h022ffd2f12d0be36022ffd2f12b0bd35022ffd2f1290bc34022ffd2f12e2fd3b),
    .INIT_50(256'h022ffd209752067a022ffd001f001b00022ffd2500001a01022ffd2f12f0bf3b),
    .INIT_51(256'h022ffd20975223ec022ffd001d0206b6022ffd2097509c07022ffd001e020628),
    .INIT_52(256'h022ffd2f62a20733022ffd2f7282071c022ffd2097536390022ffd001c01d051),
    .INIT_53(256'h022ffd01500206de022ffd01400363ec022ffd2f42e1d020022ffd2f52c09006),
    .INIT_54(256'h022ffd2f62b1dec0022ffd2f7293a3ec022ffd01700206cc022ffd016000120a),
    .INIT_55(256'h022ffd001f0223ec022ffd2294132358022ffd2f42f0de80022ffd2f52d32364),
    .INIT_56(256'h022ffd001d00ba02022ffd20975206a2022ffd001e0206a2022ffd20975206a2),
    .INIT_57(256'h022ffd001702fc0c022ffd20975206a2022ffd001c0363ec022ffd2097518fa0),
    .INIT_58(256'h022ffd001602237a022ffd037f02ff0f022ffd2f1292fe0e022ffd0310f2fd0d),
    .INIT_59(256'h022ffd001500ba02022ffd036f0206a2022ffd2f12b206a2022ffd0310f206a2),
    .INIT_5A(256'h022ffd001402fc10022ffd035f0206a2022ffd2f12d363ec022ffd0310f18ea0),
    .INIT_5B(256'h022ffd011000b105022ffd034f00b004022ffd2f12f2fe12022ffd0310f2fd11),
    .INIT_5C(256'h022ffd2f12e1ae20022ffd2f12c1ad10022ffd2f12a18c00022ffd2f1280b206),
    .INIT_5D(256'h022ffd1410003401022ffd144000b40f022ffd1410020b5f022ffd229413e3ec),
    .INIT_5E(256'h022ffd14100208fa022ffd1460020896022ffd141002237a022ffd145002f40f),
    .INIT_5F(256'h022ffd141000127b022ffd144002b6c9022ffd141002b00a022ffd14700206dc),
    .INIT_60(256'h022ffd1410009c08022ffd1460009d08022ffd1410009e08022ffd1450009f08),
    .INIT_61(256'h022ffd0b82800ce0022ffd00170206b6022ffd2500000cd0022ffd14700206b6),
    .INIT_62(256'h022ffd20a51206dc022ffd20a33206b6022ffd20a2700cf0022ffd0b929206b6),
    .INIT_63(256'h022ffd14b00223ed022ffd14a0e208a5022ffd0ba2536380022ffd01b0019201),
    .INIT_64(256'h022ffd14a0020733022ffd14b002071a022ffd14a00363ee022ffd0ba261d050),
    .INIT_65(256'h022ffd0b217206de022ffd14b00363ec022ffd14a001d020022ffd14b0009006),
    .INIT_66(256'h022ffd14b00206a2022ffd14a003a3ec022ffd2f217206cc022ffd062b001202),
    .INIT_67(256'h022ffd14b0018bc0022ffd14a000bc02022ffd14b00206a2022ffd14a00206a2),
    .INIT_68(256'h022ffd14b0009002022ffd14a00206a2022ffd14b00206a2022ffd14a00363ec),
    .INIT_69(256'h022ffd14a001fb00022ffd14b001da00022ffd14a00363da022ffd0ba270d040),
    .INIT_6A(256'h022ffd0b216323da022ffd14b001fb00022ffd14a001da20022ffd14b00323da),
    .INIT_6B(256'h022ffd0b82a1daa0022ffd00160323da022ffd2fb161fb00022ffd06b201da80),
    .INIT_6C(256'h022ffd20a511fb00022ffd20a331dac0022ffd20a27323da022ffd0b92b1fb00),
    .INIT_6D(256'h022ffd14b00323da022ffd14a0e1fb00022ffd0ba251dae0022ffd01b00323da),
    .INIT_6E(256'h022ffd14a001da80022ffd14b00323da022ffd14a001fb01022ffd0ba261da20),
    .INIT_6F(256'h022ffd0b2191fb01022ffd14b001daa0022ffd14a00323da022ffd14b001fb01),
    .INIT_70(256'h022ffd14b00323da022ffd14a001fb01022ffd2f2191dac0022ffd062b0323da),
    .INIT_71(256'h022ffd14b001da20022ffd14a00323da022ffd14b001fb02022ffd14a001da00),
    .INIT_72(256'h022ffd14b001fb02022ffd14a001da80022ffd14b00323da022ffd14a001fb02),
    .INIT_73(256'h022ffd14a00323da022ffd14b001fb02022ffd14a001daa0022ffd0ba27323da),
    .INIT_74(256'h022ffd0b2181da00022ffd14b00323da022ffd14a001fb02022ffd14b001dac0),
    .INIT_75(256'h022ffd0b82c1fb03022ffd001501dae0022ffd2fb18323da022ffd06b201fb03),
    .INIT_76(256'h022ffd20a5120896022ffd20a33206dc022ffd20a27223ec022ffd0b92d323da),
    .INIT_77(256'h022ffd14b00208b7022ffd14a0e208d4022ffd0ba25001b0022ffd01b00000a0),
    .INIT_78(256'h022ffd14a00206b6022ffd14b0000cf0022ffd14a0000bc0022ffd0ba26208e4),
    .INIT_79(256'h022ffd0b21b206b6022ffd14b0000cd0022ffd14a00206b6022ffd14b0000ce0),
    .INIT_7A(256'h022ffd14b00223ec022ffd14a00208a5022ffd2f21b206b6022ffd062b000cb0),
    .INIT_7B(256'h022ffd14b0020718022ffd14a0022008022ffd14b002077b022ffd14a00206dc),
    .INIT_7C(256'h022ffd14b00208a5022ffd14a0020137022ffd14b0020896022ffd14a00206dc),
    .INIT_7D(256'h022ffd14a0001002022ffd14b002b80f022ffd14a002b40f022ffd0ba272b20f),
    .INIT_7E(256'h022ffd0b21a206dc022ffd14b0022008022ffd14a002077b022ffd14b002074d),
    .INIT_7F(256'h022ffd0b82e2b20f02bff300140208a502bff02fb1a20137022ffd06b2020896),
    .INITP_00(256'h61d3daf741ce5d617e514b55ecd1f3f87a6348d761eec142ce7e56f4635fd75a),
    .INITP_01(256'he6e8dcf4417a426e7fe04df879f046eddf734b76d27e567d4adedf61eae0d66f),
    .INITP_02(256'h7c6cec7fe7e2d5e2fd4feae241e5f9cb717741e2f9ceea71417bea49e76bdf66),
    .INITP_03(256'h465bfce76cef76eb7b68f34e797462ebfaf77cff4f6160e27ff874f1e4cbf8f5),
    .INITP_04(256'heee3db7673feecc04fd2707a4fe14d50e57d51f9c46a70ea4969cf7a62ebdaf3),
    .INITP_05(256'h6154f5e26f79c1d17aefef4c4155d37ec742f2fbe565e2e479fcfe6aed71f5f5),
    .INITP_06(256'hd14d5ff46bd2d8dbee4d6ad07675e0c462cb6be165f669eaf162edf5fbf37d7f),
    .INITP_07(256'he1e0e142e8d16050f049d8745fdee773fe5c635df8eed865fc45c744fa4763fc),
    .INITP_08(256'h55df4cc5d8ce5ec34f405fd15a5de9f56873c76ed375dbee5c69e67543dc4745),
    .INITP_09(256'hda584d59cdc0d5c4dee94d7b5f69526642525ccd72cd6573476369dfcfdbf4e8),
    .INITP_0A(256'hd24370cee943734373f74cede9cbcce164d256e57fcad6fdddfdcf7d4a78f54e),
    .INITP_0B(256'hedfff96078da75c2f5e2787f55cedec1c1634e7b5bc7d7e04b404c6049fbc173),
    .INITP_0C(256'hecd66f4c6fd14ec64773567ec7ead56172c6eec3cbed6ffb4b406b63e649e8c0),
    .INITP_0D(256'h4666c4fdcfe7def6e747f0c2d66ae87e5f59c5f05c7ec9e75d6050e4f84c6f50),
    .INITP_0E(256'hf34de5d952eefe60c6524664c1e7d8e7c4fb45e1fbcfe7d8eac4fb43e7de59c2),
    .INITP_0F(256'h55e8f0e65979cbe8ceefd276ffc0fa406f5ae840f1dc454e40ea43e94360cc6b),
