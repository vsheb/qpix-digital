    .INIT_00(256'h00b8340d0ff20020022bf8012002ff00032c2f2066b01f0001c2d03260628000),
    .INIT_01(256'h0012000b11b2078702f20f0b01a0100100ba362f2212004900b9351420020033),
    .INIT_02(256'h032cc11f1ff1d00201d4011d0ff3205d0094082f1151d0010013002f01420778),
    .INIT_03(256'h03ac160d0ff1d01001ba00012003225601b9002066b1d0000188403261232136),
    .INIT_04(256'h02f9350b11d1d00802f8340b01c325360133002f2221d0040112011420032472),
    .INIT_05(256'h00b9351d0ff0106000b8342f1153221d022c092f0141d08202fa3601200325d5),
    .INIT_06(256'h02f80c012002074402f20d2066b2078702f30e3261f0109f00ba361f1ff2077b),
    .INIT_07(256'h00b70f2084622ffd00b60e2f2232071600b50d142002075c00b40c0d0ff2074c),
    .INIT_08(256'h0147000b1210b0000146080b0203202f0146082084b0d08000b30e2089409002),
    .INIT_09(256'h00b0020b123011ff02f70e04010010ff0147000b1223602f014308040100d001),
    .INIT_0A(256'h014006050401b200014006207751b1000140063262d19001014006040100121f),
    .INIT_0B(256'h00b4392077b09001025000030bf2f000037000207750100102f00f2262f3e029),
    .INIT_0C(256'h00b43c190012b000032c650b01f2500001d4002f03b3202f0034f00b00e0d040),
    .INIT_0D(256'h01ba002b40f0900101b9002b20f2be0f018840208e02bf7e0012003663b2b00c),
    .INIT_0E(256'h02f9352f01f0d02002f834226600900d011201010022d00103ac402b80f0300f),
    .INIT_0F(256'h022c351d00209006032c65220082203a01d2022079d0900602fa36010823603f),
    .INIT_10(256'h02f20f1d0103604600ba363265a0d08000b9351d0080900d00b8343265a09006),
    .INIT_11(256'h01b90020775090070188403664c090070194021d0202204100b43c3265a09007),
    .INIT_12(256'h00b935226602074e00b834010022073e03ecc12077b2075a01ba000504025000),
    .INIT_13(256'h003301030bf2075c000380207752074c00b20f366532075e00ba361d0402071a),
    .INIT_14(256'h02f80d1d0802076002f30c226602071a014808010022073601490e2077b20758),
    .INIT_15(256'h0142002077b20716014908030bf2071e014908207752071a0003903601720720),
    .INIT_16(256'h001302208e03e05a02f20e2011e1900101420622660010190143080100225000),
    .INIT_17(256'h01400601000200bc0140062077b200d601400605040200ce00b0022077525000),
    .INIT_18(256'h0370000900d208d102f30f2200832060004300207b50d001014006207870900d),
    .INIT_19(256'h0188400900d208f2001200250002090f00b43836663011010250000d08001080),
    .INIT_1A(256'h011201014400100003ac72250003606301ba00366671dc9301b9000d0402091f),
    .INIT_1B(256'h01c2d00b0142f00202fa360b2150100002f935013002f00102f8340150a05001),
    .INIT_1C(256'h00b9350d0081d11200b834143000311e022c6714200001e0032c940d01020bd1),
    .INIT_1D(256'h019402011010100000b438030072208002f20f143000120200ba361420032077),
    .INIT_1E(256'h03ecc1226781400001ba00141060dd4001b9003a67c3607e018840190010dd10),
    .INIT_1F(256'h00b20f2d2090122100ba362d30a2f00200b935123501400000b834102400dd20),
    .INIT_20(256'h00039001a002f03a02f80d250000100002f30c02010200b8001300090082f239),
    .INIT_21(256'h01430809c1c2f02401420014b060100101490814b060d0040149080bb1309002),
    .INIT_22(256'h00b00210ba0208dd00130309f1f200f202f20e09e1e200c801420009d1d200e1),
    .INIT_23(256'h01400613f002094801400613e002b02e01400613d00208e001400610cb0208da),
    .INIT_24(256'h02500020663200b8037000206ad208d102f30f01b002094800430001a042b02e),
    .INIT_25(256'h01b900206632b04e01884009d07200b8001200206632011000b40309c07200c2),
    .INIT_26(256'h02f83401a73320ad01120109f071d00103ac9f206630300f01ba0009e0709001),
    .INIT_27(256'h00b8340b612208e0022c960b511320a702fa360b4100d00202f93501b0109002),
    .INIT_28(256'h00b40312e600100202f20f12d502b80f00ba3610c402b40f00b935036012b20f),
    .INIT_29(256'h01ba003e6a12011e01b9001bb002200801884019a01207b501940213f0020787),
    .INIT_2A(256'h00ba36206ad207b500b93501b012078700b83401a740100003ecc125000208e0),
    .INIT_2B(256'h02f80d206672b40f02f30c2df072b20f00130020667208e000b20f2500022008),
    .INIT_2C(256'h01420020667207a30149082dd072f03201490820667010010003902de072b80f),
    .INIT_2D(256'h00130420667224bf02f20e2db0720718014200206672071c0143082dc072073c),
    .INIT_2E(256'h01400601500250000140060146c20716014006250002074a00b0022da0720752),
    .INIT_2F(256'h0370000d0102075402f30f0b014207360043000b2152073a0140060130020746),
    .INIT_30(256'h02f20d142002075002f20c0d008207460012ff14300250000250001420020718),
    .INIT_31(256'h0250001900125000037000011012071802f20f030072075c02f20e1430020746),
    .INIT_32(256'h020ce5102402074a00b117226c72073800b016141062073c0013003a6cb20758),
    .INIT_33(256'h001301090082075a02f2202d2092074002f1172d30a2500002f0161235020718),
    .INIT_34(256'h02f0182d008206ef020ce52d2090300f00b1192d30a0900100b0180601020718),
    .INIT_35(256'h00b01a14c002074000130214b002073602f22114a062500002f1192500020716),
    .INIT_36(256'h02f11b250001400e02f01a14f0003008020ce514e000900200b11b14d0020718),
    .INIT_37(256'h00b11d14c082071600b01c14d08206ef00130314e081400e02f22214f0e1400e),
    .INIT_38(256'h02f223110b92090f02f11d250000110002f01c14a08010c0020ce514b0825000),
    .INIT_39(256'h01f1ff1901101c0001d0ff3900001d00001200190e901e020250003900001f00),
    .INIT_3A(256'h014006190f62090f014006390000110301400611007010000310003e6ed20929),
    .INIT_3B(256'h01410000c0001c000140062500001d000141001100a01e000140062500001f00),
    .INIT_3C(256'h010030206f70110001400e2076a010c001400e207012500001400e206f720929),
    .INIT_3D(256'h022ffd0110001d01022ffd2500001e000250002076a01f0000b224207012090f),
    .INIT_3E(256'h022ffd1410001100022ffd14c06010a0022ffd1410020929022ffd14c0601c00),
    .INIT_3F(256'h022ffd1410001d00022ffd14c0601e00022ffd1410001f00022ffd14c062090f),
    .INIT_40(256'h022ffd1110701101022ffd3a704010c0022ffd1d10a20929022ffd2500001c00),
    .INIT_41(256'h022ffd2076d03e3c022ffd01a0003f81022ffd2500020926022ffd111302090f),
    .INIT_42(256'h022ffd0110405e40022ffd3900005f00022ffd206e303c3f022ffd0900603d7c),
    .INIT_43(256'h022ffd04a0025000022ffd3670c20929022ffd1910105c00022ffd206d505d03),
    .INIT_44(256'h022ffd1920120926022ffd2076a2090f022ffd2070101101022ffd00100010c0),
    .INIT_45(256'h022ffd2276a03cff022ffd0110d03dfd022ffd2500003e7f022ffd3670703fff),
    .INIT_46(256'h022ffd2276a05c00022ffd0115f05d00022ffd2276a05e80022ffd0112005f00),
    .INIT_47(256'h022ffd2276a01101022ffd01131010c0022ffd2276a25000022ffd0113e20929),
    .INIT_48(256'h022ffd2276a03eff022ffd0113003fff022ffd2276a20926022ffd011332090f),
    .INIT_49(256'h022ffd2276a25000022ffd0113220929022ffd2276a03cff022ffd0113103dfe),
    .INIT_4A(256'h022ffd2276a20926022ffd011342090f022ffd2276a01101022ffd01133010c0),
    .INIT_4B(256'h022ffd2276a03cff022ffd0113603dfe022ffd2276a03eff022ffd0113503fff),
    .INIT_4C(256'h022ffd2276a05c00022ffd0113805d01022ffd2276a05e00022ffd0113705f00),
    .INIT_4D(256'h022ffd2276a2f032022ffd0114101000022ffd2276a25000022ffd0113920929),
    .INIT_4E(256'h022ffd2276a3617c022ffd011430d040022ffd2276a0900f022ffd011422f01e),
    .INIT_4F(256'h022ffd2276a36177022ffd011450d080022ffd2276a3617c022ffd011440d020),
    .INIT_50(256'h022ffd2276a0d040022ffd0114736173022ffd2276a0d080022ffd011460900e),
    .INIT_51(256'h022ffd2276a0d010022ffd011493616d022ffd2276a0d020022ffd0114836170),
    .INIT_52(256'h022ffd2276a32153022ffd0114b0d004022ffd2276a0900e022ffd0114a3616a),
    .INIT_53(256'h022ffd2276a0300f022ffd0114d2b04e022ffd2276a2f033022ffd0114c09016),
    .INIT_54(256'h022ffd2276a0900d022ffd0114f22161022ffd2276a36160022ffd0114e1d00e),
    .INIT_55(256'h022ffd2276a1d049022ffd0115109006022ffd2276a36160022ffd011500d020),
    .INIT_56(256'h022ffd2276a36160022ffd011531d053022ffd2276a22161022ffd011523615a),
    .INIT_57(256'h022ffd2276a207b5022ffd01155207be022ffd2276a20716022ffd011542075a),
    .INIT_58(256'h022ffd2276a208d1022ffd0115720716022ffd2276a20746022ffd0115622008),
    .INIT_59(256'h022ffd2276a20787022ffd0115901000022ffd2276a208e0022ffd011582011e),
    .INIT_5A(256'h022ffd2d10601080022ffd207712b10e022ffd2276a22008022ffd0115a207b5),
    .INIT_5B(256'h022ffd3676d2217a022ffd0d02001040022ffd0900d2b20e022ffd250002217a),
    .INIT_5C(256'h022ffd36771208d1022ffd0d0102217a022ffd0900d01020022ffd250002b40e),
    .INIT_5D(256'h022ffd25000208d1022ffd030602217a022ffd0900001010022ffd250002b80e),
    .INIT_5E(256'h022ffd00100221f3022ffd250002f01e022ffd0309f01008022ffd090002b80f),
    .INIT_5F(256'h022ffd2d10001001022ffd041002b20f022ffd207782b40f022ffd03160208d1),
    .INIT_60(256'h022ffd207750b237022ffd2071819801022ffd2073a0982f022ffd207402f01e),
    .INIT_61(256'h022ffd00100208f2022ffd250002090f022ffd2071601102022ffd206ef010a0),
    .INIT_62(256'h022ffd2d1002fd0d022ffd041002fc0c022ffd2077503f07022ffd0319f2091f),
    .INIT_63(256'h022ffd0b0320bd0d022ffd207180bc0c022ffd2073a2ff0f022ffd2075a2fe0e),
    .INIT_64(256'h022ffd206ef01100022ffd2077801020022ffd327b10bf0f022ffd1d0010be0e),
    .INIT_65(256'h022ffd2073a0d001022ffd2075a0b001022ffd2500020929022ffd207162090f),
    .INIT_66(256'h022ffd20716208e6022ffd206ef2219e022ffd0100222017022ffd207183619b),
    .INIT_67(256'h022ffd207751d000022ffd0319f0b016022ffd001002094c022ffd25000208fe),
    .INIT_68(256'h022ffd010001f000022ffd250000b018022ffd2d1001f000022ffd041000b017),
    .INIT_69(256'h022ffd2075a1f000022ffd2d1030b01a022ffd0b1321f000022ffd2079d0b019),
    .INIT_6A(256'h022ffd1d0011f000022ffd0b0320b01c022ffd207181f000022ffd2073a0b01b),
    .INIT_6B(256'h022ffd207160b032022ffd206ef361ba022ffd010401f000022ffd327b10b01d),
    .INIT_6C(256'h022ffd2071611001022ffd206ef0b03a022ffd0102032512022ffd250001d002),
    .INIT_6D(256'h022ffd327bc1d001022ffd1d0000b032022ffd20778208e0022ffd250002f03a),
    .INIT_6E(256'h022ffd250000d001022ffd207180b001022ffd2071c22008022ffd20752324bf),
    .INIT_6F(256'h022ffd207500b016022ffd2075a321f0022ffd227b91d800022ffd2074630935),
    .INIT_70(256'h022ffd207160b018022ffd206f02f035022ffd0bc020b017022ffd207182f034),
    .INIT_71(256'h022ffd207460b01a022ffd207582f03b022ffd207800b019022ffd2078c2f036),
    .INIT_72(256'h022ffd207160b01c022ffd206f02f03d022ffd0bc3a0b01b022ffd207182f03c),
    .INIT_73(256'h022ffd207182092c022ffd207402f03f022ffd2074e0b01d022ffd250002f03e),
    .INIT_74(256'h022ffd206f00b016022ffd0bc062094c022ffd20722208fe022ffd20722208e6),
    .INIT_75(256'h022ffd206f00b135022ffd0bc040b017022ffd206f01c010022ffd0bc050b134),
    .INIT_76(256'h022ffd207381e010022ffd2075c0b136022ffd208230b018022ffd207161e010),
    .INIT_77(256'h022ffd3a7e20b01a022ffd0d5041e010022ffd095020b13b022ffd207180b019),
    .INIT_78(256'h022ffd09d1d0b13d022ffd09c1c0b01b022ffd227f91e010022ffd208350b13c),
    .INIT_79(256'h022ffd14b061e010022ffd0bb020b13e022ffd09f1f0b01c022ffd09e1e1e010),
    .INIT_7A(256'h022ffd13e0036202022ffd13d001e010022ffd10cb00b13f022ffd14b060b01d),
    .INIT_7B(256'h022ffd2fd35221cf022ffd2fe36321f0022ffd2ff3b1d800022ffd13f0019801),
    .INIT_7C(256'h022ffd0bc360b002022ffd206f02f01f022ffd0bc3b01004022ffd2fc3420af7),
    .INIT_7D(256'h022ffd0bc34321f9022ffd206f01d002022ffd0bc350b032022ffd206f02f013),
    .INIT_7E(256'h022ffd207381d001022ffd2073a0b032022ffd20716207c6022ffd206f020716),
    .INIT_7F(256'h022ffd2083501004022ffd3a80132536022ffd0d5041d002022ffd2071832536),
    .INITP_00(256'ha00025b46949d9293339cdd95063b425679a81ba6b8e9382904da4198ef7e99f),
    .INITP_01(256'hf742a2dd7677a863acb28a9bbb741c9d2c7c7ddea0243b260d66bd98a394192d),
    .INITP_02(256'h3d2b383081571f129987859ee4e22d909380b9830295473a242eaf147e35baa6),
    .INITP_03(256'h23269491d4a9a43bbf2ffd0190b17747814a656b225e388b9f2d11df59dc0937),
    .INITP_04(256'h1f49c94f5b81f23715a182194ac4d786248d8c02b4aa770bb50f0ca439e3603a),
    .INITP_05(256'he16ab130332f338288ef27302f19a2ad5652b13c27a63e479927a18492e83fb3),
    .INITP_06(256'h9caa956348f4cca719bc70ef4d462db210f2f759d71734316acf6bd8ee548f74),
    .INITP_07(256'hf95df753e74b7d535ff97e9c151234863a203d2eac90006a3a14b942f2d07dc4),
    .INITP_08(256'h5bd3d6c35f77dd59dbd2657fc36351efe3f9defc5cc8f2c8616ff9fb7777f6f7),
    .INITP_09(256'hc465c579c565477d5674d65e5fd7515adb49d545c54c5b48d642dbd4d543c5d1),
    .INITP_0A(256'hd6f4d665cd62ccf2cdfccdfbc277cde7416bd5705c75c4f2ddf3de625f64d8f8),
    .INITP_0B(256'h6359e1c0f1617f41f06b4fedcce0d7f35bfbc678eb67c4f550774ce8cc6e5466),
    .INITP_0C(256'h74d77bfd46e0685b40797ec2f7f2634c635fddedf4db6dccfdf754fc68d7cbec),
    .INITP_0D(256'h7675cf6aeb43cbe670c4e16d497d7dfb5c6ec972da7a42cc786cd3696861644e),
    .INITP_0E(256'h666a52cd46705743697ee8e5e8f955db54e5f3ebd2606441ee606ce35467f946),
    .INITP_0F(256'h40f0e744cdc2d167fd766aeee86f766bd743747a57504f627058d27ae954f74f),
