    .INIT_00(256'h00b8340150001f0103ec7a0146c2ff0001ba002500001f0001b9002da0728000),
    .INIT_01(256'h0003800d0102202a00b20f0b0142202a00ba360b2152800000b935013002df02),
    .INIT_02(256'h02f30c142002df020148080d00801f0001490e143002202a003301142002202a),
    .INIT_03(256'h014908190013201d014908011011d00400039003007206c302f80d1430028000),
    .INIT_04(256'h02f20e10240325420142062260f1d00101430814106325ba0142003a6131d002),
    .INIT_05(256'h014006090081d0000140062d2093209100b0132d30a1d00200130212350206c0),
    .INIT_06(256'h02f30f2d0081d0820043002d209324dc0140062d30a1d0100140060601032282),
    .INIT_07(256'h00120014c002800000b43814b002df0202500014a0601f010370002500032225),
    .INIT_08(256'h03ac2b250002202a01ba0014f002202a01b90014e002202a01884014d002202a),
    .INIT_09(256'h02fa3614c082202a02f93514d082202a02f83414e082202a01120114f0e2202a),
    .INIT_0A(256'h00b834110b9206c6022c202500001060032c4d14a082202a01c2d014b082202a),
    .INIT_0B(256'h00b438190112069402f20f390002068c00ba36190e9206d200b935390000109f),
    .INIT_0C(256'h01ba00190f6010c001b9003900022ffc018840110072065e0194023e635206a4),
    .INIT_0D(256'h00ba3600c00208d500b935250002500000b8341100a208b703ec7a2500001101),
    .INIT_0E(256'h02f80d2063f03cff02f30c206b203dfe0013002064903eff00b20f2063f03fff),
    .INIT_0F(256'h0142000110020033014908250002079f014908206b22500000039020649208e5),
    .INIT_10(256'h001303141000110002f20e14c0620037014200141000110001430814c0601010),
    .INIT_11(256'h014006141002089501400614c062500001400614100208ce00b01314c0601014),
    .INIT_12(256'h037000111072003702f30f3a64c011000043001d10a010140140062500020033),
    .INIT_13(256'h018840206b52500000120001a00208ce00b40325000010140250001113001100),
    .INIT_14(256'h011201011040110003ac58390000101801ba002062b2003301b900090062089b),
    .INIT_15(256'h022c4f04a00208ce02fa36366540101802f935191010110002f8342061d20037),
    .INIT_16(256'h02f20f192010101c00ba36206b22003300b93520649208a500b8340010025000),
    .INIT_17(256'h01b900226b2011000188400110d0101c019402250002003700b4033664f01100),
    .INIT_18(256'h00b935226b203fff00b8340115f208d503ec7a226b22500001ba0001120208ce),
    .INIT_19(256'h02f30c226b205f000013000113103cff00b20f226b203dfe00ba360113e03eff),
    .INIT_1A(256'h014908226b2208e50149080113005c00000390226b205d0102f80d0113305e00),
    .INIT_1B(256'h02f20e226b2010100142000113220033014308226b22079f0142000113125000),
    .INIT_1C(256'h014006226b201014014006011340110000b013226b2200620013040113301100),
    .INIT_1D(256'h02f30f226b2200330043000113620895014006226b22500001400601135208ce),
    .INIT_1E(256'h02f20c226b2011000012ff0113820062025000226b2011000370000113701014),
    .INIT_1F(256'h037000226b22089b02f20f011412500002f20e226b2208ce02f20d0113901014),
    .INIT_20(256'h022ffc226b220062022ffc0114301100022ffc226b2010180250000114220033),
    .INIT_21(256'h022ffc226b225000022ffc01145208ce022ffc226b201018022ffc0114401100),
    .INIT_22(256'h022ffc226b201100022ffc011470101c022ffc226b220033022ffc01146208a5),
    .INIT_23(256'h022ffc226b2208ce022ffc0114901100022ffc226b20101c022ffc0114820062),
    .INIT_24(256'h022ffc226b22f01e022ffc0114b2f032022ffc226b201000022ffc0114a25000),
    .INIT_25(256'h022ffc226b209012022ffc0114d320c4022ffc226b20d008022ffc0114c09011),
    .INIT_26(256'h022ffc226b2320a9022ffc0114f1d004022ffc226b2320a0022ffc0114e1d008),
    .INIT_27(256'h022ffc226b2320bb022ffc011511d001022ffc226b2320b2022ffc011501d002),
    .INIT_28(256'h022ffc226b20d040022ffc011530900f022ffc226b22f001022ffc0115201000),
    .INIT_29(256'h022ffc226b20d080022ffc0115536112022ffc226b20d020022ffc0115436112),
    .INIT_2A(256'h022ffc226b20900f022ffc011572f001022ffc226b201001022ffc011563610c),
    .INIT_2B(256'h022ffc226b236112022ffc011590d004022ffc226b236112022ffc011580d008),
    .INIT_2C(256'h022ffc2d1062f001022ffc206b901002022ffc226b23610c022ffc0115a0d010),
    .INIT_2D(256'h022ffc366b50d020022ffc0d02036112022ffc0900d0d040022ffc2500009010),
    .INIT_2E(256'h022ffc366b901003022ffc0d0103610c022ffc0900d0d080022ffc2500036112),
    .INIT_2F(256'h022ffc2500036112022ffc030600d008022ffc0900009010022ffc250002f001),
    .INIT_30(256'h022ffc090133610c022ffc250000d010022ffc0309f36112022ffc090000d004),
    .INIT_31(256'h022ffc031600d040022ffc0010036107022ffc250000d080022ffc030070900e),
    .INIT_32(256'h022ffc206880d010022ffc2d100360ff022ffc041000d020022ffc206c036103),
    .INIT_33(256'h022ffc20637320d7022ffc206bd0d004022ffc206600900e022ffc20682360fb),
    .INIT_34(256'h022ffc0319f0300f022ffc001002b04e022ffc250002f033022ffc2065e09016),
    .INIT_35(256'h022ffc206a20900d022ffc2d100220ea022ffc04100360e9022ffc206bd1d00e),
    .INIT_36(256'h022ffc1d0011d049022ffc0b03209006022ffc20660360e9022ffc206820d020),
    .INIT_37(256'h022ffc2065e360e9022ffc206371d053022ffc206c0220ea022ffc326fc360de),
    .INIT_38(256'h022ffc2066001300022ffc206820b202022ffc206a22065e022ffc25000206a2),
    .INIT_39(256'h022ffc25000360e4022ffc2065e1c320022ffc2063711301022ffc010022071c),
    .INIT_3A(256'h022ffc041002065e022ffc206bd2068e022ffc0319f2200a022ffc0010020713),
    .INIT_3B(256'h022ffc206e81d002022ffc010000b002022ffc2500020047022ffc2d1002003e),
    .INIT_3C(256'h022ffc206821d003022ffc206a20b002022ffc2d10320050022ffc0b132320f6),
    .INIT_3D(256'h022ffc326fc01000022ffc1d0012085b022ffc0b03220059022ffc20660320f6),
    .INIT_3E(256'h022ffc250002b10e022ffc2065e2200a022ffc2063720713022ffc01040206d2),
    .INIT_3F(256'h022ffc250002b20e022ffc2065e22110022ffc2063701080022ffc0102020700),
    .INIT_40(256'h022ffc2b04f2b40e022ffc2b08f22110022ffc2b20f01040022ffc2b40f20700),
    .INIT_41(256'h022ffc2d01020887022ffc0102022110022ffc2d01001020022ffc0104020700),
    .INIT_42(256'h022ffc2d01022110022ffc0100401010022ffc2d01020700022ffc010082b80e),
    .INIT_43(256'h022ffc2d01001008022ffc0108020700022ffc2b10f0b001022ffc2b80f20887),
    .INIT_44(256'h022ffc206c020047022ffc250002003e022ffc2d010221ed022ffc010102f01e),
    .INIT_45(256'h022ffc2066420050022ffc2069a3211c022ffc3271a1d002022ffc1d0000b002),
    .INIT_46(256'h022ffc2271720059022ffc2068e3211c022ffc250001d003022ffc206600b002),
    .INIT_47(256'h022ffc00c302f01e022ffc2066001001022ffc2069820700022ffc206a20b001),
    .INIT_48(256'h022ffc206cb0b001022ffc206d70b237022ffc2065e19801022ffc206380982f),
    .INIT_49(256'h022ffc0bc3a32137022ffc206601d001022ffc2068e3212c022ffc206a01d000),
    .INIT_4A(256'h022ffc00c3032155022ffc250001d003022ffc2065e32145022ffc206381d002),
    .INIT_4B(256'h022ffc20660208e2022ffc20688208b7022ffc2069601102022ffc2fc13010a0),
    .INIT_4C(256'h022ffc0bc062fe0e022ffc20b7a2fd0d022ffc2066a2fc0c022ffc2066a03f07),
    .INIT_4D(256'h022ffc0bc042079f022ffc2063822167022ffc0bc05208e8022ffc206382ff0f),
    .INIT_4E(256'h022ffc206a401102022ffc20784010a0022ffc2065e2079f022ffc2063820855),
    .INIT_4F(256'h022ffc0d5042fc0c022ffc0950203f07022ffc20660208e2022ffc20680208b7),
    .INIT_50(256'h022ffc09c1c208eb022ffc2275a2ff0f022ffc207962fe0e022ffc3a7432fd0d),
    .INIT_51(256'h022ffc0bb132079f022ffc09f1f20855022ffc09e1e2079f022ffc09d1d2216a),
    .INIT_52(256'h022ffc13d0001102022ffc10cb0010a0022ffc14b062079f022ffc14b0620855),
    .INIT_53(256'h022ffc2fe362fc0c022ffc2ff3b03f07022ffc13f00208e2022ffc13e00208b7),
    .INIT_54(256'h022ffc20638208ee022ffc0bc3b2ff0f022ffc2fc342fe0e022ffc2fd352fd0d),
    .INIT_55(256'h022ffc206382079f022ffc0bc3520855022ffc206382079f022ffc0bc362216d),
    .INIT_56(256'h022ffc206822079f022ffc2065e20855022ffc206382079f022ffc0bc3420855),
    .INIT_57(256'h022ffc3a762208e2022ffc0d504208b7022ffc2066001102022ffc20680010a0),
    .INIT_58(256'h022ffc0bd352fe0e022ffc0bc342fd0d022ffc227782fc0c022ffc2079603f07),
    .INIT_59(256'h022ffc01b00207cd022ffc01a0422170022ffc0bf3b208f1022ffc0be362ff0f),
    .INIT_5A(256'h022ffc205ed2093c022ffc09f07207d4022ffc205ed22172022ffc205f52093c),
    .INIT_5B(256'h022ffc205ed22172022ffc09d072093c022ffc205ed207de022ffc09e0722172),
    .INIT_5C(256'h022ffc206381d000022ffc00cd00b016022ffc206382093c022ffc09c07207ea),
    .INIT_5D(256'h022ffc206381f000022ffc00cf00b018022ffc206381f000022ffc00ce00b017),
    .INIT_5E(256'h022ffc206601f000022ffc206940b01a022ffc206821f000022ffc2065e0b019),
    .INIT_5F(256'h022ffc14c001f000022ffc0d5040b01c022ffc01c001f000022ffc2066a0b01b),
    .INIT_60(256'h022ffc250000b032022ffc2065e36199022ffc206381f000022ffc11c010b01d),
    .INIT_61(256'h022ffc2b80c11001022ffc206600b03a022ffc206a2325ba022ffc206a41d002),
    .INIT_62(256'h022ffc2b02c0b002022ffc2063820076022ffc09c0c2006d022ffc2b03c2f03a),
    .INIT_63(256'h022ffc09c0c0b002022ffc2b01c2007f022ffc2063832193022ffc09c0c1d002),
    .INIT_64(256'h022ffc2063820700022ffc09c0c20088022ffc2b00c32193022ffc206381d003),
    .INIT_65(256'h022ffc206ac32542022ffc206ac1d001022ffc250000b032022ffc2065e2085b),
    .INIT_66(256'h022ffc206ac0b016022ffc206ac321e8022ffc206ac1d800022ffc206ac2200a),
    .INIT_67(256'h022ffc2bec90b018022ffc250002f035022ffc206ac0b017022ffc206ac2f034),
    .INIT_68(256'h022ffc209280b01a022ffc2b08e2f03b022ffc2b1bb0b019022ffc2b21a2f036),
    .INIT_69(256'h022ffc207b80b01c022ffc01c002f03d022ffc250000b01b022ffc208b32f03c),
    .INIT_6A(256'h022ffc250000b001022ffc207b82f03f022ffc01c100b01d022ffc250002f03e),
    .INIT_6B(256'h022ffc01c0d321b8022ffc250001d001022ffc207b8321b4022ffc01c071d000),
    .INIT_6C(256'h022ffc207b8321c0022ffc01c011d003022ffc25000321bc022ffc207b81d002),
    .INIT_6D(256'h022ffc25000221c3022ffc207b82093c022ffc01c04207cd022ffc25000208e8),
    .INIT_6E(256'h022ffc208c0221c3022ffc01f002093c022ffc01e00207d4022ffc01d00208eb),
    .INIT_6F(256'h022ffc207c7221c3022ffc208b72093c022ffc01100207de022ffc01080208ee),
    .INIT_70(256'h022ffc2b63b0b016022ffc2b00a2093c022ffc2b389207ea022ffc25000208f1),
    .INIT_71(256'h022ffc2b2090b135022ffc250000b017022ffc209281c010022ffc2b08e0b134),
    .INIT_72(256'h022ffc209281e010022ffc2b08e0b136022ffc2b37b0b018022ffc2b00a1e010),
    .INIT_73(256'h022ffc2b62a0b01a022ffc2b6491e010022ffc207b50b13b022ffc250000b019),
    .INIT_74(256'h022ffc250000b13d022ffc209280b01b022ffc2b08e1e010022ffc2b5bb0b13c),
    .INIT_75(256'h022ffc207b51e010022ffc2079f0b13e022ffc208550b01c022ffc2079f1e010),
    .INIT_76(256'h022ffc2b08e361ff022ffc2b5bb1e010022ffc2b62a0b13f022ffc2b6490b01d),
    .INIT_77(256'h022ffc208550b001022ffc2079f321e8022ffc250001d800022ffc2092819801),
    .INIT_78(256'h022ffc207b5321b8022ffc2079f1d001022ffc20855321b4022ffc2079f1d000),
    .INIT_79(256'h022ffc2b08e321c0022ffc2b5bb1d003022ffc2b62a321bc022ffc2b6491d002),
    .INIT_7A(256'h022ffc2085501004022ffc2079f20aa0022ffc250002f013022ffc209280b001),
    .INIT_7B(256'h022ffc208550b032022ffc2079f2f013022ffc208550b001022ffc2079f2f01f),
    .INIT_7C(256'h022ffc2b62a20724022ffc2b6492065e022ffc207b5321f3022ffc2079f1d002),
    .INIT_7D(256'h022ffc250001d002022ffc20928321fc022ffc2b08e1d001022ffc2b5bb0b032),
    .INIT_7E(256'h022ffc2bdfb2200a022ffc2b10a206d2022ffc2b64901004022ffc207b2321fc),
    .INIT_7F(256'h022ffc2b10a0b03a022ffc2b6c92200a022ffc209282d003022ffc2b08e01004),
    .INITP_00(256'h008a4c75cf0b868916bc1caefeb884a118200f5473bc350d0f36a6911845a99e),
    .INITP_01(256'hac06b98f634e2dae339eb6ccb21d8f0f82f01db78ffb490651e27d03480e22a0),
    .INITP_02(256'ha90b0526e3ba23077979d1f594ddb88397a3a0f662ed8533a494270e95dc84a2),
    .INITP_03(256'h7b4ff64e5c10e5c1f9b62f852385bb1e68b69b348e202141efb7b2b08f035e9a),
    .INITP_04(256'h57d1d3cd5b50dfcbc0db5fdf51ded944cecbd1ddd4d4d951da505750d8cd57eb),
    .INITP_05(256'h5353754041467f53cd4af85acee8c1d14c5f4cc44bc45a40d44cd25653cc5f44),
    .INITP_06(256'hf1c65357694d6afbf85673e2e0d9c6735b7666e1fe5865557c5ecbe7eecec2ee),
    .INITP_07(256'h5d7e59555e78d36dc96658f0616cc9ff5a4048cd6c7de041d96043d9747dedc1),
    .INITP_08(256'h6ef4e16a427457f4ecf663e844c466d575e8cbd3e056fb5aea4ef8ebd65dc2c1),
    .INITP_09(256'h40fa6bf0e052e7c655cfda4ad4dbebff6b6dfa5e6c57efc74b6377e35342fd5c),
    .INITP_0A(256'hfa41ff6dfbffdeccded6dedc4840cbf77fd358fc68e9cbd3f4e0c1d46de440f7),
    .INITP_0B(256'h61d444fff3e474e7516d51744276ce715f4f4a45d2f15fd16e4ecb7ff7cb65df),
    .INITP_0C(256'hc6c5fa7579f2f361f9e146fb5ce5e244e8f8db7970dbede95ff0607a46f451fc),
    .INITP_0D(256'heecb63fcf75c657b5c4fd058de4bc546ded250ca43d5d3c45ac4484bc2d27a54),
    .INITP_0E(256'hd2d1c0de4fcb7a4750da5949cc414addf855c6cd50de5ef443c9435bfd70c955),
    .INITP_0F(256'hcffcdf5347474c5ad4c7c1d470c840c4d75cd2ddd14a4c4a5fc5f6d84ac25341),
