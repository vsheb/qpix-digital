library IEEE;
use IEEE.STD_LOGIC_1164.all;

package QpixPkg is

   -- Define some enums for making directional connections
   constant RT : integer := 0;
   constant DN : integer := 1;
   constant LT : integer := 2;
   constant UP : integer := 3;
   
end QpixPkg;

package body QpixPkg is

end package body QpixPkg;
