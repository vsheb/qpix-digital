    localparam [35:0] init1FB = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init1FC = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init1FD = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init1FE = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init1FF = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init200 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init201 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init202 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init203 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init204 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init205 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init206 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init207 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init208 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init209 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init20A = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init20B = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init20C = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init20D = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init20E = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init20F = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init210 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init211 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init212 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init213 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init214 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init215 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init216 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init217 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init218 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init219 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init21A = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init21B = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init21C = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init21D = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init21E = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init21F = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init220 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init221 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init222 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init223 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init224 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init225 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init226 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init227 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init228 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init229 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init22A = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init22B = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init22C = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init22D = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init22E = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init22F = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init230 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init231 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init232 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init233 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init234 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init235 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init236 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init237 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init238 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init239 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init23A = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init23B = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init23C = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init23D = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init23E = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init23F = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init240 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init241 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init242 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init243 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init244 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init245 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init246 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init247 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init248 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init249 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init24A = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init24B = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init24C = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init24D = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init24E = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init24F = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init250 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init251 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init252 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init253 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init254 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init255 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init256 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init257 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init258 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init259 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init25A = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init25B = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init25C = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init25D = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init25E = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init25F = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init260 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init261 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init262 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init263 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init264 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init265 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init266 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init267 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init268 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init269 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init26A = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init26B = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init26C = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init26D = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init26E = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init26F = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init270 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init271 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init272 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init273 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init274 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init275 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init276 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init277 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init278 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init279 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init27A = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init27B = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init27C = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init27D = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init27E = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init27F = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init280 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init281 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init282 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init283 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init284 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init285 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init286 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init287 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init288 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init289 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init28A = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init28B = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init28C = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init28D = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init28E = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init28F = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
