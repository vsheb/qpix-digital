    .INIT_00(256'h022bfc2b02c20528022bfc204c62200a022bfc09c0c204ee022bfc2b03c204f2),
    .INIT_01(256'h022bfc09c0c2051c022bfc2b01c25000022bfc204c6204ec022bfc09c0c20520),
    .INIT_02(256'h022bfc204c6204ee022bfc09c0c2052a022bfc2b00c2050c022bfc204c620510),
    .INIT_03(256'h022bfc2053a2051c022bfc2053a20526022bfc250002051c022bfc204ec25000),
    .INIT_04(256'h022bfc2053a2052e022bfc2053a25000022bfc2053a204ee022bfc2053a20532),
    .INIT_05(256'h022bfc0b032204ee022bfc2500020520022bfc2053a2050e022bfc2053a20512),
    .INIT_06(256'h022bfc20528204ee022bfc2051020530022bfc3661e20516022bfc1d00025000),
    .INIT_07(256'h022bfc20510204ec022bfc25000204c5022bfc204ec0300f022bfc2052e09001),
    .INIT_08(256'h022bfc25000204ee022bfc204ec20516022bfc2050c2050c022bfc2052225000),
    .INIT_09(256'h022bfc205141400e022bfc3662b1400e022bfc1d00003008022bfc0b03209002),
    .INIT_0A(256'h022bfc2500025000022bfc204ec204ec022bfc20512204c5022bfc205261400e),
    .INIT_0B(256'h022bfc204ec01f00022bfc20510207be022bfc2051001100022bfc20514010c0),
    .INIT_0C(256'h022bfc204ee207ec022bfc2050c01c00022bfc2052a01d00022bfc205fc01e02),
    .INIT_0D(256'h022bfc14106207be022bfc1410601103022bfc1410601000022bfc0b11325000),
    .INIT_0E(256'h022bfc204c501c00022bfc0401001d00022bfc0b00f01e00022bfc1410601f00),
    .INIT_0F(256'h022bfc204c501100022bfc0b00d010c0022bfc204c525000022bfc0b00e207ec),
    .INIT_10(256'h022bfc2052201d01022bfc204ec01e00022bfc204c501f00022bfc0b00c207be),
    .INIT_11(256'h022bfc204c5010a0022bfc0100025000022bfc204ee207ec022bfc2050c01c00),
    .INIT_12(256'h022bfc0b01201e00022bfc1410601f00022bfc14106207be022bfc0b11301100),
    .INIT_13(256'h022bfc204c525000022bfc0b011207ec022bfc204c501c00022bfc0401001d00),
    .INIT_14(256'h022bfc2500003d7c022bfc204ec03e3c022bfc204c503f81022bfc0b010207dc),
    .INIT_15(256'h022bfc0bc1605d02022bfc3469205e40022bfc1dcff05f00022bfc0bc1703c3f),
    .INIT_16(256'h022bfc1dcff207dc022bfc0bc1925000022bfc34698207ec022bfc1dcff05c00),
    .INIT_17(256'h022bfc3469803cff022bfc1dcff03dfd022bfc0bc1803e7f022bfc3469203fff),
    .INIT_18(256'h022bfc0bc1a05c00022bfc3469205d00022bfc1dcff05e80022bfc0bc1b05f00),
    .INIT_19(256'h022bfc1dcff01101022bfc0bc1d010c0022bfc3469825000022bfc1dcff207ec),
    .INIT_1A(256'h022bfc3469803fff022bfc1dcff207dc022bfc0bc1c25000022bfc34692207be),
    .INIT_1B(256'h022bfc32676207ec022bfc1dd0003cff022bfc0bd2003dfe022bfc2500003eff),
    .INIT_1C(256'h022bfc2069e01010022bfc0bc1620266022bfc20692206aa022bfc0bc1725000),
    .INIT_1D(256'h022bfc1dd0001010022bfc0bd2101100022bfc206a42026a022bfc0bc2001100),
    .INIT_1E(256'h022bfc0bc1820266022bfc20692207a0022bfc0bc1925000022bfc3267f207d5),
    .INIT_1F(256'h022bfc0bd2201100022bfc206a42026a022bfc0bc2101100022bfc2069e01014),
    .INIT_20(256'h022bfc20692207a6022bfc0bc1b25000022bfc32688207d5022bfc1dd0001014),
    .INIT_21(256'h022bfc206a42026a022bfc0bc2201100022bfc2069e01018022bfc0bc1a20266),
    .INIT_22(256'h022bfc0bc1d25000022bfc32691207d5022bfc1dd0001018022bfc0bd2301100),
    .INIT_23(256'h022bfc0bc2301100022bfc2069e0101c022bfc0bc1c20266022bfc20692207b0),
    .INIT_24(256'h022bfc20512207d5022bfc2053801100022bfc250000101c022bfc206a42026a),
    .INIT_25(256'h022bfc2500003eff022bfc204ee03fff022bfc204c6207dc022bfc204ee25000),
    .INIT_26(256'h022bfc204c605e00022bfc204ee05f00022bfc2053203cff022bfc2050e03dfe),
    .INIT_27(256'h022bfc2053225000022bfc2050e207ec022bfc2500005c00022bfc204ec05d01),
    .INIT_28(256'h022bfc2500001100022bfc204ee01010022bfc204c620266022bfc204ee206aa),
    .INIT_29(256'h022bfc204c6207d5022bfc204ee01010022bfc2053601100022bfc2052220295),
    .INIT_2A(256'h022bfc2b21a01014022bfc2bec920266022bfc25000207a0022bfc204ec25000),
    .INIT_2B(256'h022bfc2007301014022bfc2082f01100022bfc2b08e20295022bfc2b1bb01100),
    .INIT_2C(256'h022bfc2500020266022bfc206c3207a6022bfc01c0025000022bfc25000207d5),
    .INIT_2D(256'h022bfc01c0701100022bfc2500020295022bfc206c301100022bfc01c1001018),
    .INIT_2E(256'h022bfc206c3207b0022bfc01c0d25000022bfc25000207d5022bfc206c301018),
    .INIT_2F(256'h022bfc2500020295022bfc206c301100022bfc01c010101c022bfc2500020266),
    .INIT_30(256'h022bfc01d0025000022bfc25000207d5022bfc206c301100022bfc01c040101c),
    .INIT_31(256'h022bfc0108001200022bfc207c73632d022bfc01f001d001022bfc01e000b01e),
    .INIT_32(256'h022bfc250002f816022bfc206d220843022bfc207be0b517022bfc011000b416),
    .INIT_33(256'h022bfc2b08e0b519022bfc2b63b0b418022bfc2b00a04210022bfc2b3892f917),
    .INIT_34(256'h022bfc2b00a04210022bfc2b2092f919022bfc250002f818022bfc2082f20843),
    .INIT_35(256'h022bfc250002f81a022bfc2082f20843022bfc2b08e0b51b022bfc2b37b0b41a),
    .INIT_36(256'h022bfc2b5bb0b51d022bfc2b62a0b41c022bfc2b64904210022bfc206c02f91b),
    .INIT_37(256'h022bfc206aa04210022bfc250002f91d022bfc2082f2f81c022bfc2b08e20843),
    .INIT_38(256'h022bfc2b6492f21e022bfc206c001202022bfc206aa322ef022bfc207600d202),
    .INIT_39(256'h022bfc2082f0b032022bfc2b08e20624022bfc2b5bb20617022bfc2b62a2062c),
    .INIT_3A(256'h022bfc206aa32398022bfc207601d002022bfc206aa32372022bfc250001d001),
    .INIT_3B(256'h022bfc2b64901204022bfc206c02236e022bfc206aa05020022bfc207602054b),
    .INIT_3C(256'h022bfc2082f0b117022bfc2b08e0b016022bfc2b5bb208a5022bfc2b62a2f21e),
    .INIT_3D(256'h022bfc206aa1f1ff022bfc207601d0ff022bfc206aa2f115022bfc250002f014),
    .INIT_3E(256'h022bfc206aa2f014022bfc207600b119022bfc206aa0b018022bfc2076034490),
    .INIT_3F(256'h022bfc2b5bb34490022bfc2b62a1f1ff022bfc2b6491d0ff022bfc206c02f115),
    .INIT_40(256'h022bfc206bd2f115022bfc250002f014022bfc2082f0b11b022bfc2b08e0b01a),
    .INIT_41(256'h022bfc2b08e0b01c022bfc2bdfb34490022bfc2b10a1f1ff022bfc2b6491d0ff),
    .INIT_42(256'h022bfc2bebb1d0ff022bfc2b10a2f115022bfc2b6c92f014022bfc2082f0b11d),
    .INIT_43(256'h022bfc206aa1d000022bfc250000b032022bfc2082f34490022bfc2b08e1f1ff),
    .INIT_44(256'h022bfc206aa3231a022bfc207541d000022bfc207e30b013022bfc01ccc36321),
    .INIT_45(256'h022bfc2bdfb3231e022bfc2b10a1d002022bfc2b6493231c022bfc206bd1d001),
    .INIT_46(256'h022bfc2b10a22321022bfc2b6c920804022bfc2082f32320022bfc2b08e1d003),
    .INIT_47(256'h022bfc2500022321022bfc2082f20819022bfc2b08e22321022bfc2bebb2080e),
    .INIT_48(256'h022bfc2075420654022bfc207e320617022bfc01cd82062c022bfc206aa20824),
    .INIT_49(256'h022bfc2075432372022bfc207e31d001022bfc01ccc0b032022bfc206aa20624),
    .INIT_4A(256'h022bfc2b10a030df022bfc2b6492054b022bfc206bd32398022bfc206aa1d002),
    .INIT_4B(256'h022bfc2b6c920510022bfc2082f3633a022bfc2b08e1d008022bfc2bdfb2236e),
    .INIT_4C(256'h022bfc2082f205fc022bfc2b08e204ec022bfc2bebb20510022bfc2b10a2052e),
    .INIT_4D(256'h022bfc207e32054b022bfc01ce432372022bfc206aa1d001022bfc250000b032),
    .INIT_4E(256'h022bfc207e336347022bfc01cd81d010022bfc206aa2236e022bfc2075405020),
    .INIT_4F(256'h022bfc207e3204ec022bfc01ccc2053a022bfc206aa20534022bfc207542050c),
    .INIT_50(256'h022bfc2b64932372022bfc206bd1d001022bfc206aa0b032022bfc20754205fc),
    .INIT_51(256'h022bfc2082f1d020022bfc2b08e2236e022bfc2bdfb05020022bfc2b10a2054b),
    .INIT_52(256'h022bfc2b08e2053a022bfc2bebb20534022bfc2b10a2050c022bfc2b6c936354),
    .INIT_53(256'h022bfc2b22a1d001022bfc2b1c90b032022bfc25000205fc022bfc2082f204ec),
    .INIT_54(256'h022bfc250002236e022bfc2082f030df022bfc2b08e2054b022bfc2b47b32372),
    .INIT_55(256'h022bfc2b08e20534022bfc2b57b2050c022bfc2b22a36361022bfc2b4891d040),
    .INIT_56(256'h022bfc2b66a0b032022bfc2b5c9205fc022bfc25000204ec022bfc2082f2053a),
    .INIT_57(256'h022bfc25000030df022bfc2082f2054b022bfc2b08e32372022bfc2b6bb1d001),
    .INIT_58(256'h022bfc2b08e2052e022bfc2b7bb3602a022bfc2b66a1d080022bfc2b6c92236e),
    .INIT_59(256'h022bfc20760205fc022bfc206aa204ec022bfc2500020524022bfc2082f20528),
    .INIT_5A(256'h022bfc207be2054b022bfc0110132372022bfc010801d001022bfc206aa0b032),
    .INIT_5B(256'h022bfc01c0e01008022bfc206aa20554022bfc250002236e022bfc206cc030df),
    .INIT_5C(256'h022bfc206b12027a022bfc206aa20271022bfc207542200a022bfc207e320560),
    .INIT_5D(256'h022bfc207e320283022bfc01c1e3237c022bfc206aa1d002022bfc250000b002),
    .INIT_5E(256'h022bfc01c0e2028c022bfc206b13237c022bfc206aa1d003022bfc207540b002),
    .INIT_5F(256'h022bfc206b101000022bfc206aa20554022bfc2075401060022bfc207e320766),
    .INIT_60(256'h022bfc207e32b20f022bfc01c2e2b40f022bfc206aa2d003022bfc250002f032),
    .INIT_61(256'h022bfc01c1e2d010022bfc206b101040022bfc206aa2b04f022bfc207542b08f),
    .INIT_62(256'h022bfc206b12d010022bfc206aa01008022bfc207542d010022bfc207e301020),
    .INIT_63(256'h022bfc206aa2b10f022bfc207542b80f022bfc207e32d010022bfc01c0e01004),
    .INIT_64(256'h022bfc1d0022d010022bfc0b00201010022bfc250002d010022bfc206b101080),
    .INIT_65(256'h022bfc1d0042200a022bfc3279b2058e022bfc1d00320560022bfc3279901000),
    .INIT_66(256'h022bfc207750b01e022bfc2279e2200a022bfc2076e2d003022bfc3279d01002),
    .INIT_67(256'h022bfc250000d004022bfc0b00209002022bfc207813640c022bfc2279e1d004),
    .INIT_68(256'h022bfc2075401f0a022bfc207e32047f022bfc01c0e20459022bfc206aa323f0),
    .INIT_69(256'h022bfc01c1a20439022bfc206aa0120b022bfc25000011b3022bfc206aa01e40),
    .INIT_6A(256'h022bfc01c0e2dd08022bfc206aa2de09022bfc207542df0a022bfc207e309d07),
    .INIT_6B(256'h022bfc25000363b1022bfc206aa1cf20022bfc20754363b1022bfc207e31ce10),
    .INIT_6C(256'h022bfc20754223a7022bfc207e313f00022bfc01c2611e01022bfc206aa223b4),
    .INIT_6D(256'h022bfc207542f115022bfc207e32f014022bfc01c1a0b117022bfc206aa0b016),
    .INIT_6E(256'h022bfc2075420441022bfc207e3323c0022bfc01c0e1f1ff022bfc206aa1d0ff),
    .INIT_6F(256'h022bfc2b4192f220022bfc2b00a14200022bfc250000d0ff022bfc206aa01200),
    .INIT_70(256'h022bfc2b2592f115022bfc2b00a2f014022bfc2d1080b119022bfc2d0080b018),
    .INIT_71(256'h022bfc2b00a20441022bfc25000323cc022bfc2d1081f1ff022bfc2d0081d0ff),
    .INIT_72(256'h022bfc2de082f221022bfc2dd0814200022bfc2dc080d0ff022bfc2b28901200),
    .INIT_73(256'h022bfc2b2892f115022bfc2b00a2f014022bfc250000b11b022bfc2df080b01a),
    .INIT_74(256'h022bfc09f0820441022bfc09e08323d8022bfc09d081f1ff022bfc09c081d0ff),
    .INIT_75(256'h022bfc2dc082f222022bfc2d00914200022bfc2d10a0d0ff022bfc2500001200),
    .INIT_76(256'h022bfc250002f014022bfc2df0801200022bfc2de080b11d022bfc2dd080b01c),
    .INIT_77(256'h022bfc09d08323e5022bfc09c081f1ff022bfc2d0091d0ff022bfc2d10a2f115),
    .INIT_78(256'h022bfc0105014200022bfc250000d0ff022bfc09f0801200022bfc09e0820441),
    .INIT_79(256'h022bfc2dc0820624022bfc2d0092066d022bfc2d10a2061f022bfc011022f223),
    .INIT_7A(256'h022bfc250000b122022bfc207ce04010022bfc206cc0b121022bfc250000b020),
    .INIT_7B(256'h022bfc206aa323f3022bfc2500004010022bfc206d20b123022bfc207c704010),
    .INIT_7C(256'h022bfc207fb2054b022bfc207a0223f5022bfc2500005040022bfc207fb2054b),
    .INIT_7D(256'h022bfc250002f03b022bfc207fb0b00e022bfc207a620554022bfc25000030bf),
    .INIT_7E(256'h022bfc01020202a0022bfc2500036408022bfc207fb19001022bfc207b00b01f),
    .INIT_7F(256'h022bfc0be0e3240502d0030bf0f1d0020010ff207be0b00202bff001100202a9),
    .INITP_00(256'h6f77dd64f6edd3d16172f3fb7973f371ff7ef04ad35d535e5dc856df40c4515f),
    .INITP_01(256'hdce4d2e7cf79e8e6f9f0fbc7d768fd61546b64f27c4ffa7b614dc672fc447070),
    .INITP_02(256'h5dd5745855e156d9e0dada71f6c8d060d279cf79ede6f9c9d779d768e359cc7b),
    .INITP_03(256'h51d9f3597158e1d17bd0d9e9df6bd7fbd1fc477f5e55e757dd795056e9d25bf0),
    .INITP_04(256'heee8f54dd45be36d7fdf56d170e677d9685e6dd1fdd77c4bd972d8ea5b7acefd),
    .INITP_05(256'h74ff6bf6f4e1fd7ce974ff69f67e7afd5fc567c5e77ef04ad25bfc78725bd9d2),
    .INITP_06(256'h4a6d54f5e2cdf262e05160ed53636551e5cf53e661efe75ad6d2ea5659fdff6d),
    .INITP_07(256'he0c6e7f7c1eb43e041794f75cae07acafbe3d560caff456b48e460c3f5f84fe7),
    .INITP_08(256'h635170dcedc341fde4e378dcc3e747655cffc5e6d875db4862677be74c754b61),
    .INITP_09(256'hc8fdc976d2675b6e43f7dfff4a6a42f8dfdefcfa6bfec9d9feda7b43f043f653),
    .INITP_0A(256'he545e27e6dd479ce6ee8fc48ef52e1437df3fdce6a4ef742d5fc747cfddc4bf2),
    .INITP_0B(256'h4948f1c565c35af34f77d9fcc84be4c86448ef68e7cdcc4b6fcdf4c265d5f641),
    .INITP_0C(256'h78f371ccfe49e7725a7f55ebd6eae0c5d0f751e5d6ccef446242d6ead6e5dbfc),
    .INITP_0D(256'h69ccfdc5724ae95ff4c4e347e3d664d7e459eb526149f948ecc4fbd0efcbef4c),
    .INITP_0E(256'he64446f47542efe6cfccf2714b60675ad1d8fc416df6495bd07a615c4cd8ed40),
    .INITP_0F(256'hcf47856f68634d7878cfea64407ae0404af0f1427bc5f0f343d5fa455bfd4768),
