    .INIT_00(256'h022ffd0be3611001022ffd0bd350b03a022ffd0bc3422008022ffd2281720787),
    .INIT_01(256'h022ffd206ad0b017022ffd01b001d000022ffd01a040b016022ffd0bf3b2f03a),
    .INIT_02(256'h022ffd09e070b019022ffd206631f000022ffd09f070b018022ffd206631f000),
    .INIT_03(256'h022ffd09c070b01b022ffd206631f000022ffd09d070b01a022ffd206631f000),
    .INIT_04(256'h022ffd00ce00b01d022ffd206f01f000022ffd00cd00b01c022ffd206f01f000),
    .INIT_05(256'h022ffd207160b032022ffd206f0208e0022ffd00cf036017022ffd206f01f000),
    .INIT_06(256'h022ffd2072232512022ffd207181d002022ffd2074c324bf022ffd2073a1d001),
    .INIT_07(256'h022ffd11c010bd10022ffd14c002f01e022ffd0d50401001022ffd01c0022008),
    .INIT_08(256'h022ffd2075c13e00022ffd2500011d01022ffd207160bf12022ffd206f00be11),
    .INIT_09(256'h022ffd2b03c03f01022ffd2b80c2fe11022ffd207182fd10022ffd2075a13f00),
    .INIT_0A(256'h022ffd09c0c03007022ffd2b02c0b00f022ffd206f020bec022ffd09c0c2ff12),
    .INIT_0B(256'h022ffd206f00be0e022ffd09c0c0307e022ffd2b01c0b03b022ffd206f02f00f),
    .INIT_0C(256'h022ffd2071620935022ffd206f03624e022ffd09c0c1c0e0022ffd2b00c03e7e),
    .INIT_0D(256'h022ffd207640b017022ffd207641d000022ffd207640b016022ffd250002094c),
    .INIT_0E(256'h022ffd207640b019022ffd207641f000022ffd207640b018022ffd207641f000),
    .INIT_0F(256'h022ffd1d0000b01b022ffd0b0321f000022ffd250000b01a022ffd207641f000),
    .INIT_10(256'h022ffd207580b01d022ffd207521f000022ffd2073a0b01c022ffd368451f000),
    .INIT_11(256'h022ffd2074c20796022ffd2073a2224e022ffd2500036247022ffd207161f000),
    .INIT_12(256'h022ffd0b03201004022ffd25000207c6022ffd2071620716022ffd20736207b5),
    .INIT_13(256'h022ffd207502b20f022ffd2073e208e0022ffd3685222008022ffd1d00020787),
    .INIT_14(256'h022ffd2073e20787022ffd2500001002022ffd207162b80f022ffd2073c2b40f),
    .INIT_15(256'h022ffd208232f032022ffd2071601000022ffd2073a22008022ffd2073a207b5),
    .INIT_16(256'h022ffd0b11309017022ffd2071832289022ffd207360d004022ffd207540900e),
    .INIT_17(256'h022ffd1410609019022ffd141062f008022ffd1410609018022ffd141062f007),
    .INIT_18(256'h022ffd0b00e0901b022ffd206ef2f00a022ffd040100901a022ffd0b00f2f009),
    .INIT_19(256'h022ffd0b00c2b04e022ffd206ef2f033022ffd0b00d09016022ffd206ef2f00b),
    .INIT_1A(256'h022ffd2073609002022ffd2074c3626f022ffd207161d00a022ffd206ef0300f),
    .INIT_1B(256'h022ffd0b1131d00e022ffd206ef22430022ffd010003242f022ffd207180d002),
    .INIT_1C(256'h022ffd040103627c022ffd0b0121d00b022ffd141062242f022ffd1410636272),
    .INIT_1D(256'h022ffd0b01020758022ffd206ef2dc01022ffd0b01103c0f022ffd206ef0bc07),
    .INIT_1E(256'h022ffd0bc1722003022ffd2500020716022ffd20716206f0022ffd206ef20718),
    .INIT_1F(256'h022ffd1dcff2244c022ffd0bc162075e022ffd348b936280022ffd1dcff1d00d),
    .INIT_20(256'h022ffd348b92243c022ffd1dcff2073c022ffd0bc1936284022ffd348bf1d00f),
    .INIT_21(256'h022ffd0bc1b32455022ffd348bf0d008022ffd1dcff32455022ffd0bc181d00c),
    .INIT_22(256'h022ffd1dcff3642f022ffd0bc1a0d020022ffd348b90900d022ffd1dcff2242d),
    .INIT_23(256'h022ffd348b909002022ffd1dcff36293022ffd0bc1d1d04f022ffd348bf09006),
    .INIT_24(256'h022ffd250001d053022ffd348bf22430022ffd1dcff3242f022ffd0bc1c0d002),
    .INIT_25(256'h022ffd0bc17207be022ffd3289d20716022ffd1dd002075a022ffd0bd203629a),
    .INIT_26(256'h022ffd0bc20362b1022ffd208c51d052022ffd0bc162242e022ffd208b9207cd),
    .INIT_27(256'h022ffd328a61d020022ffd1dd0009006022ffd0bd212076d022ffd208cb20758),
    .INIT_28(256'h022ffd208c509006022ffd0bc182076d022ffd208b920718022ffd0bc193642d),
    .INIT_29(256'h022ffd1dd002076d022ffd0bd2220722022ffd208cb3642d022ffd0bc211d030),
    .INIT_2A(256'h022ffd0bc1a2d001022ffd208b93a42d022ffd0bc1b206e3022ffd328af09006),
    .INIT_2B(256'h022ffd0bd2320716022ffd208cb2076a022ffd0bc2220701022ffd208c500100),
    .INIT_2C(256'h022ffd208b92075e022ffd0bc1d362b5022ffd328b81d055022ffd1dd0022003),
    .INIT_2D(256'h022ffd208cb2073c022ffd0bc23362b9022ffd208c51d044022ffd0bc1c2244c),
    .INIT_2E(256'h022ffd2071820750022ffd2073c362e0022ffd207621d04e022ffd250002243c),
    .INIT_2F(256'h022ffd207383642d022ffd250001d020022ffd2071809006022ffd206f02076d),
    .INIT_30(256'h022ffd207163a42d022ffd206f020706022ffd207180120a022ffd2075c20718),
    .INIT_31(256'h022ffd207182fd0b022ffd2075c2fc0a022ffd207382fb09022ffd250002fa08),
    .INIT_32(256'h022ffd2074c3a42d022ffd2500020706022ffd2071801201022ffd206f02fe33),
    .INIT_33(256'h022ffd2071614a06022ffd206f014a06022ffd2071814a06022ffd2076014a06),
    .INIT_34(256'h022ffd2b1bb0be0b022ffd2b00a0bd0a022ffd2b0090bc09022ffd250000bb08),
    .INIT_35(256'h022ffd208e9206dc022ffd01c00206dc022ffd20944206dc022ffd2b08e0bf33),
    .INIT_36(256'h022ffd208e92fc09022ffd01c102fb08022ffd250002fa07022ffd20059206dc),
    .INIT_37(256'h022ffd2500022466022ffd208e92ff33022ffd01c072fe0b022ffd250002fd0a),
    .INIT_38(256'h022ffd01c012076d022ffd250002075c022ffd208e936350022ffd01c0d1d054),
    .INIT_39(256'h022ffd208e920718022ffd01c043642d022ffd250001d020022ffd208e909006),
    .INIT_3A(256'h022ffd01f002fa08022ffd01e003a42d022ffd01d0020706022ffd250000120a),
    .INIT_3B(256'h022ffd2090f2fe33022ffd011002fd0b022ffd010802fc0a022ffd209182fb09),
    .INIT_3C(256'h022ffd2b00a3a42d022ffd2b3893a42d022ffd2500020706022ffd208f801201),
    .INIT_3D(256'h022ffd2500014a06022ffd2094414a06022ffd2b08e14a06022ffd2b63b14a06),
    .INIT_3E(256'h022ffd2b08e0bc09022ffd2b37b0bb08022ffd2b00a0ba07022ffd2b1c92fa07),
    .INIT_3F(256'h022ffd2b62a206dc022ffd2b6490bf33022ffd250000be0b022ffd209440bd0a),
    .INIT_40(256'h022ffd250002fa07022ffd20944206dc022ffd2b08e206dc022ffd2b5bb206dc),
    .INIT_41(256'h022ffd2b08e2fe0b022ffd2bdcb2fd0a022ffd2b10a2fc09022ffd2b6492fb08),
    .INIT_42(256'h022ffd2bebb1df0c022ffd2b10a2fb3f022ffd2b6c92fa3e022ffd209442ff33),
    .INIT_43(256'h022ffd2b00a2242d022ffd2500032310022ffd209440df08022ffd2b08e32330),
    .INIT_44(256'h022ffd2b00a206d5022ffd2d1083642d022ffd2d00818fa0022ffd2b4190ba02),
    .INIT_45(256'h022ffd250002fc0c022ffd2d108206d5022ffd2d008206d5022ffd2b259206d5),
    .INIT_46(256'h022ffd2dd0820af7022ffd2dc082ff0f022ffd2b2892fe0e022ffd2b00a2fd0d),
    .INIT_47(256'h022ffd2b00a0bf12022ffd250000be11022ffd2df080bd10022ffd2de0820716),
    .INIT_48(256'h022ffd09e08206f0022ffd09d0800cf0022ffd09c0820722022ffd2b2892073a),
    .INIT_49(256'h022ffd2091f206f0022ffd208f200cd0022ffd25000206f0022ffd09f0800ce0),
    .INIT_4A(256'h022ffd2500020701022ffd208f8206f7022ffd20918206f7022ffd250000bc3f),
    .INIT_4B(256'h022ffd0bf0f2242d022ffd2090f206f0022ffd011000bc3e022ffd010202076a),
    .INIT_4C(256'h022ffd2092918ea0022ffd0bc0c0ba02022ffd0bd0d206d5022ffd0be0e206d5),
    .INIT_4D(256'h022ffd208fe2fc10022ffd208e6206d5022ffd2092c206d5022ffd250003642d),
    .INIT_4E(256'h022ffd2092c20bec022ffd2500003e03022ffd2093b2fe12022ffd250002fd11),
    .INIT_4F(256'h022ffd208f20bd0e022ffd2090f0be0d022ffd011010bf0c022ffd0108020716),
    .INIT_50(256'h022ffd25000206f0022ffd2090400cd0022ffd208e3206f0022ffd208f80bc0f),
    .INIT_51(256'h022ffd25000206f0022ffd3694400cf0022ffd0d008206f0022ffd0900e00ce0),
    .INIT_52(256'h022ffd2500020701022ffd32948206f7022ffd0d002206f7022ffd0900e0bc3f),
    .INIT_53(256'h022ffd2f1172242d022ffd2f116206f0022ffd011000bc3e022ffd370012076a),
    .INIT_54(256'h022ffd2f11b0d004022ffd2f11a09002022ffd2f1193636e022ffd2f1181d058),
    .INIT_55(256'h022ffd2b6c909006022ffd010a22076d022ffd2f11d20764022ffd2f11c3e36e),
    .INIT_56(256'h022ffd2096201208022ffd1100120718022ffd2b00b3642d022ffd2b00a1d020),
    .INIT_57(256'h022ffd3695a2fa34022ffd1d0ff20716022ffd209c13a42d022ffd2096720706),
    .INIT_58(256'h022ffd09d080bc34022ffd09c082fd3b022ffd250002fc36022ffd370002fb35),
    .INIT_59(256'h022ffd1d0d001a01022ffd250000bf3b022ffd09f080be36022ffd09e080bd35),
    .INIT_5A(256'h022ffd001f009c07022ffd3299220663022ffd1d0d1206ad022ffd3297d01b00),
    .INIT_5B(256'h022ffd001d0363d1022ffd209b01d051022ffd001e02242d022ffd209b0206f0),
    .INIT_5C(256'h022ffd011001d020022ffd209b009006022ffd001c02076d022ffd209b020756),
    .INIT_5D(256'h022ffd2f12e20706022ffd2f12c0120a022ffd2f12a20718022ffd2f1283642d),
    .INIT_5E(256'h022ffd2f12f2fc0a022ffd2f12d2fb09022ffd2f12b2fa08022ffd2f1293a42d),
    .INIT_5F(256'h022ffd001e020706022ffd209b001201022ffd001f02fe33022ffd250002fd0b),
    .INIT_60(256'h022ffd001c014a06022ffd209b014a06022ffd001d014a06022ffd209b03a42d),
    .INIT_61(256'h022ffd2f52c0bd0a022ffd2f62a0bc09022ffd2f7280bb08022ffd209b014a06),
    .INIT_62(256'h022ffd01600206dc022ffd01500206dc022ffd014000bf33022ffd2f42e0be0b),
    .INIT_63(256'h022ffd2f52d2fb08022ffd2f62b2fa07022ffd2f729206dc022ffd01700206dc),
    .INIT_64(256'h022ffd209b02ff33022ffd001f02fe0b022ffd2297c2fd0a022ffd2f42f2fc09),
    .INIT_65(256'h022ffd209b032399022ffd001d00df08022ffd209b0323a5022ffd001e01df0c),
    .INIT_66(256'h022ffd0310f3642d022ffd0017018fa0022ffd209b00ba02022ffd001c02242d),
    .INIT_67(256'h022ffd0310f206d5022ffd00160206d5022ffd037f0206d5022ffd2f129206d5),
    .INIT_68(256'h022ffd0310f2ff0f022ffd001502fe0e022ffd036f02fd0d022ffd2f12b2fc0c),
    .INIT_69(256'h022ffd0310f0ba02022ffd00140206d5022ffd035f0206d5022ffd2f12d223bb),
    .INIT_6A(256'h022ffd2f128206d5022ffd01100206d5022ffd034f03642d022ffd2f12f18ea0),
    .INIT_6B(256'h022ffd2297c0b004022ffd2f12e2fe12022ffd2f12c2fd11022ffd2f12a2fc10),
    .INIT_6C(256'h022ffd145001ad10022ffd1410018c00022ffd144000b206022ffd141000b105),
    .INIT_6D(256'h022ffd147000b40f022ffd1410020bec022ffd146003e42d022ffd141001ae20),
    .INIT_6E(256'h022ffd14500208d1022ffd14100223bb022ffd144002f40f022ffd1410003407),
    .INIT_6F(256'h022ffd147002b6c9022ffd141002b00a022ffd1460020716022ffd1410020935),
    .INIT_70(256'h022ffd0b92909d08022ffd0b82809e08022ffd0017009f08022ffd250000125d),
    .INIT_71(256'h022ffd01b00206f0022ffd20a8c00cd0022ffd20a6e206f0022ffd20a6209c08),
    .INIT_72(256'h022ffd0ba26206f0022ffd14b0000cf0022ffd14a0e206f0022ffd0ba2500ce0),
    .INIT_73(256'h022ffd14b00208e0022ffd14a00363c1022ffd14b0019201022ffd14a0020716),
    .INIT_74(256'h022ffd062b020754022ffd0b2173642f022ffd14b001d050022ffd14a002242e),
    .INIT_75(256'h022ffd14a003642d022ffd14b001d020022ffd14a0009006022ffd2f2172076d),
    .INIT_76(256'h022ffd14a003a42d022ffd14b0020706022ffd14a0001202022ffd14b0020718),
    .INIT_77(256'h022ffd0ba270bc02022ffd14b00206d5022ffd14a00206d5022ffd14b00206d5),
    .INIT_78(256'h022ffd14b00206d5022ffd14a00206d5022ffd14b003642d022ffd14a0018bc0),
    .INIT_79(256'h022ffd06b201da00022ffd0b2163641b022ffd14b000d040022ffd14a0009002),
    .INIT_7A(256'h022ffd0b92b1fb00022ffd0b82a1da20022ffd001603241b022ffd2fb161fb00),
    .INIT_7B(256'h022ffd01b003241b022ffd20a8c1fb00022ffd20a6e1da80022ffd20a623241b),
    .INIT_7C(256'h022ffd0ba261dac0022ffd14b003241b022ffd14a0e1fb00022ffd0ba251daa0),
    .INIT_7D(256'h022ffd14b001fb00022ffd14a001dae0022ffd14b003241b022ffd14a001fb00),
    .INIT_7E(256'h022ffd062b03241b022ffd0b2191fb01022ffd14b001da20022ffd14a003241b),
    .INIT_7F(256'h022ffd14a001daa002bff314b003241b02bff014a001fb01022ffd2f2191da80),
    .INITP_00(256'hc24276fecfd462565cfd57e0d9e0dbe0d65d765df75d575dcfdafef35a4ee16f),
    .INITP_01(256'hcaf0e4e36ce3efe368f0ebfa43f14ccc765b59e6d75d7f50cffa59e46e6fcb78),
    .INITP_02(256'h756ff6e84ec0c4f75cdc5341db6c5b5ce2c7dec1f2e4dfc06a55f858eae54c48),
    .INITP_03(256'hd67b71507eeadcfdfc716062effdf97ac1606ec25379c96e71fa6afee97de2ef),
    .INITP_04(256'h65724152e4d463e96ce6ed4cfa7a4776f75c73f6d3fe70d4e766cd787ccee4f0),
    .INITP_05(256'h4af4d06ecd5278f255625e61ea78ec74d3d4e3db60f760e96e4ccdfc5264e2e7),
    .INITP_06(256'hf2c7667d45e1f3d4d1e4d4e449d3597a50e84af7f7634b74d1e2ca74ceee4a7c),
    .INITP_07(256'hd1fbfe48666a5dff655376d256f263d372d8d772f5594665dd60f4ccff63cfe7),
    .INITP_08(256'h53f546fae0c2d25073f2d1d1cbeed462556344fad174dac2eee9f875f3d4f170),
    .INITP_09(256'h49764f4de7ece6f54b55737a7df05a5cfb62d079e3dee175fcdae95efc73decb),
    .INITP_0A(256'h6ec569cb4e5acd5951c0c350cd4043595a51d07ae3ddf440e9fd725de9fcdcc1),
    .INITP_0B(256'hfeccfafecedfd6c2c75a5659d2576149efd7654161c54348c5f0c9efe64cf27b),
    .INITP_0C(256'he859eb5ff4c25d7ac36e417f5cfeffce79f35a4566e1d75c646fd8cde7cd7953),
    .INITP_0D(256'h78f94b75d671e1f665f1cef2d765e7e4eb54cac3454070d07b464f57f84653d1),
    .INITP_0E(256'hf3e7c4e759e2c06fd8755dc6c0df7d5cf1d8e648746051744d4441ccf2c84767),
    .INITP_0F(256'h45d9f7524a46ea4c7e4e6f5dfb6f47fb4ad0c5c77ed3d1c57c40e2dbe7c4fbcf),
