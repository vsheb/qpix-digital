    .INIT_00(256'h0013032200820020014206207632ff000142000108201f000149082f01f28000),
    .INIT_01(256'h0013013261f2074d02f20e1d008010010142083261f200490143081d00220033),
    .INIT_02(256'h02f30f366111d0020043001d0203205d0140063261f1d00100b0021d0102073e),
    .INIT_03(256'h02f20c010021d0100012ff2074132265025000050401d0000370002073b32145),
    .INIT_04(256'h0370002073b1d00802f20f36618324f102f20e1d0401d00402f20d226253242c),
    .INIT_05(256'h00b117226250106000b016010023222c001300207411d082025000030bf32590),
    .INIT_06(256'h02f220030bf2070a02f1172073b2074d02f016360170109f020c321d08020741),
    .INIT_07(256'h020c322012d22ffd00b11922625206dc00b01801002207220013012074120712),
    .INIT_08(256'h001302207410b00002f221050403202f02f1192073b0d08002f018208a509002),
    .INIT_09(256'h02f01a22008011ff020c322077b010ff00b11b2074d3602f00b01a010000d001),
    .INIT_0A(256'h00b01c250001b200001303366281b10002f2220d0801900102f11b0900d0121f),
    .INIT_0B(256'h02f11d250000900102f01c3662c2f000020c320d0400100100b11d0900d3e029),
    .INIT_0C(256'h01d0ff0bf052b0000012000be0425000025000015093202f02f223014d00d040),
    .INIT_0D(256'h0140062263a09001014006326382be0f0310001ff322bf7e01f1ff1dedb2b00c),
    .INIT_0E(256'h0140060b2150d020014100013000900d0140060150a2d001014006014400300f),
    .INIT_0F(256'h01400e143000900601400e142002203a01400e0d010090060141000b0143603f),
    .INIT_10(256'h022ffd0300736046025000143000d08000b224142000900d0100300d00809006),
    .INIT_11(256'h022ffd1410609007022ffd3a64909007022ffd1900122041022ffd0110109007),
    .INIT_12(256'h022ffd2d30a20714022ffd1235020704022ffd1024020720022ffd2264525000),
    .INIT_13(256'h022ffd2500020722022ffd0201020712022ffd0900820724022ffd2d209206e0),
    .INIT_14(256'h022ffd14b0620726022ffd14b06206e0022ffd0bb13206fc022ffd01a002071e),
    .INIT_15(256'h022ffd09f1f206dc022ffd09e1e206e4022ffd09d1d206e0022ffd09c1c206e6),
    .INIT_16(256'h022ffd13e003e05a022ffd13d0019001022ffd10cb001019022ffd10ba025000),
    .INIT_17(256'h022ffd2067a200dc022ffd01b00200f6022ffd01a04200ee022ffd13f0025000),
    .INIT_18(256'h022ffd09d0720896022ffd2062832060022ffd09c070d001022ffd206280900d),
    .INIT_19(256'h022ffd09f07208b7022ffd20628208d4022ffd09e0701101022ffd2062801080),
    .INIT_1A(256'h022ffd0b51101000022ffd0b41036063022ffd01b011dc93022ffd01aeb208e4),
    .INIT_1B(256'h022ffd12d502f002022ffd10c4001000022ffd036012f001022ffd0b61205001),
    .INIT_1C(256'h022ffd1bb001d102022ffd19a010311e022ffd13f00001e0022ffd12e6020b46),
    .INIT_1D(256'h022ffd01b011d104022ffd01aec32082022ffd250001d110022ffd3e66e32080),
    .INIT_1E(256'h022ffd2df071d116022ffd2062c32089022ffd250001d112022ffd2067a32087),
    .INIT_1F(256'h022ffd2dd0722017022ffd2062c3208d022ffd2de071d100022ffd2062c3208d),
    .INIT_20(256'h022ffd2db0701220022ffd2062c001d0022ffd2dc07320a1022ffd2062c01200),
    .INIT_21(256'h022ffd0146c01203022ffd250002208d022ffd2da07320a1022ffd2062c1d190),
    .INIT_22(256'h022ffd0b0141d190022ffd0b21501204022ffd01300001d0022ffd01500320a1),
    .INIT_23(256'h022ffd0d00836094022ffd143000dd10022ffd1420001000022ffd0d010320a1),
    .INIT_24(256'h022ffd0110114000022ffd030070dd20022ffd1430014000022ffd142000dd40),
    .INIT_25(256'h022ffd226941d112022ffd141063209b022ffd3a6981d110022ffd190012f002),
    .INIT_26(256'h022ffd2d20901222022ffd2d30a3209f022ffd123501d116022ffd102403209d),
    .INIT_27(256'h022ffd2d20901226022ffd2d30a320a1022ffd0601001223022ffd09008320a1),
    .INIT_28(256'h022ffd14b0001000022ffd14a06200d8022ffd250002f239022ffd2d008320a1),
    .INIT_29(256'h022ffd14f0001001022ffd14e000d004022ffd14d0009002022ffd14c002f03a),
    .INIT_2A(256'h022ffd190e9208a2022ffd3900020101022ffd110b9200e8022ffd250002f024),
    .INIT_2B(256'h022ffd110072090d022ffd3e6b32b02e022ffd19011208a5022ffd390002089f),
    .INIT_2C(256'h022ffd1100a200d8022ffd2500020896022ffd190f62090d022ffd390002b02e),
    .INIT_2D(256'h022ffd206c72b04e022ffd206bd200d8022ffd00c002011f022ffd25000200e2),
    .INIT_2E(256'h022ffd20730320cd022ffd206c71d001022ffd206bd0300f022ffd2073009001),
    .INIT_2F(256'h022ffd14100208a5022ffd14c06320c7022ffd011000d002022ffd2500009002),
    .INIT_30(256'h022ffd1410001002022ffd14c062b80f022ffd141002b40f022ffd14c062b20f),
    .INIT_31(256'h022ffd1d10a2012d022ffd2500022008022ffd141002077b022ffd14c062074d),
    .INIT_32(256'h022ffd250002077b022ffd111302074d022ffd1110701000022ffd3a6ca208a5),
    .INIT_33(256'h022ffd206a92b40f022ffd090062b20f022ffd20733208a5022ffd01a0022008),
    .INIT_34(256'h022ffd1910120769022ffd206a22f032022ffd0110401001022ffd390002b80f),
    .INIT_35(256'h022ffd206c72247a022ffd00100206de022ffd04a00206e2022ffd366d220702),
    .INIT_36(256'h022ffd2500025000022ffd366cd206dc022ffd1920120710022ffd2073020718),
    .INIT_37(256'h022ffd227302071a022ffd01120206fc022ffd2273020700022ffd0110d2070c),
    .INIT_38(256'h022ffd2273020716022ffd0113e2070c022ffd2273025000022ffd0115f206de),
    .INIT_39(256'h022ffd2273025000022ffd01133206de022ffd2273020722022ffd011312070c),
    .INIT_3A(256'h022ffd2273020710022ffd01131206fe022ffd2273020702022ffd011302071e),
    .INIT_3B(256'h022ffd2273020720022ffd0113320706022ffd2273025000022ffd01132206de),
    .INIT_3C(256'h022ffd22730206b5022ffd011350300f022ffd2273009001022ffd01134206de),
    .INIT_3D(256'h022ffd2273020706022ffd01137206fc022ffd2273025000022ffd01136206dc),
    .INIT_3E(256'h022ffd227301400e022ffd0113903008022ffd2273009002022ffd01138206de),
    .INIT_3F(256'h022ffd22730206dc022ffd01142206b5022ffd227301400e022ffd011411400e),
    .INIT_40(256'h022ffd22730208d4022ffd0114401100022ffd22730010c0022ffd0114325000),
    .INIT_41(256'h022ffd2273001c00022ffd0114601d01022ffd2273001e00022ffd0114501f00),
    .INIT_42(256'h022ffd22730208d4022ffd0114801100022ffd22730010a0022ffd01147208ee),
    .INIT_43(256'h022ffd2273001c00022ffd0114a01d00022ffd2273001e00022ffd0114901f00),
    .INIT_44(256'h022ffd22730208d4022ffd0114c01101022ffd22730010c0022ffd0114b208ee),
    .INIT_45(256'h022ffd2273003d7c022ffd0114e03e3c022ffd2273003f81022ffd0114d208eb),
    .INIT_46(256'h022ffd2273005d03022ffd0115005e40022ffd2273005f00022ffd0114f03c3f),
    .INIT_47(256'h022ffd22730010c0022ffd0115225000022ffd22730208ee022ffd0115105c00),
    .INIT_48(256'h022ffd2273003fff022ffd01154208eb022ffd22730208d4022ffd0115301101),
    .INIT_49(256'h022ffd2273005f00022ffd0115603cff022ffd2273003dfd022ffd0115503e7f),
    .INIT_4A(256'h022ffd22730208ee022ffd0115805c00022ffd2273005d00022ffd0115705e80),
    .INIT_4B(256'h022ffd22730208d4022ffd0115a01101022ffd22730010c0022ffd0115925000),
    .INIT_4C(256'h022ffd0900d03dfe022ffd2500003eff022ffd2d10603fff022ffd20737208eb),
    .INIT_4D(256'h022ffd0900d010c0022ffd2500025000022ffd36733208ee022ffd0d02003cff),
    .INIT_4E(256'h022ffd0900003fff022ffd25000208eb022ffd36737208d4022ffd0d01001101),
    .INIT_4F(256'h022ffd0309f05f00022ffd0900003cff022ffd2500003dfe022ffd0306003eff),
    .INIT_50(256'h022ffd2073e208ee022ffd0316005c00022ffd0010005d01022ffd2500005e00),
    .INIT_51(256'h022ffd207002f01e022ffd207062f032022ffd2d10001000022ffd0410025000),
    .INIT_52(256'h022ffd206dc0d020022ffd206b53618b022ffd2073b0d040022ffd206de0900f),
    .INIT_53(256'h022ffd2073b0900e022ffd0319f36186022ffd001000d080022ffd250003618b),
    .INIT_54(256'h022ffd207003617f022ffd207200d040022ffd2d10036182022ffd041000d080),
    .INIT_55(256'h022ffd3277736179022ffd1d0010d010022ffd0b0323617c022ffd206de0d020),
    .INIT_56(256'h022ffd250000901b022ffd206dc32162022ffd206b50d004022ffd2073e0900e),
    .INIT_57(256'h022ffd010021d0e0022ffd206de030f0022ffd207002b04e022ffd207202f00b),
    .INIT_58(256'h022ffd001000d020022ffd250000900d022ffd206dc22170022ffd206b53616f),
    .INIT_59(256'h022ffd2d10036169022ffd041001d049022ffd2073b09006022ffd0319f3616f),
    .INIT_5A(256'h022ffd0b13220720022ffd207633616f022ffd010001d053022ffd2500022170),
    .INIT_5B(256'h022ffd206de22008022ffd207002077b022ffd2072020784022ffd2d103206dc),
    .INIT_5C(256'h022ffd010402012d022ffd3277720896022ffd1d001206dc022ffd0b0322070c),
    .INIT_5D(256'h022ffd010202077b022ffd250002074d022ffd206dc01000022ffd206b5208a5),
    .INIT_5E(256'h022ffd2073e22189022ffd2500001080022ffd206dc2b10e022ffd206b522008),
    .INIT_5F(256'h022ffd206e22b40e022ffd2071822189022ffd3278201040022ffd1d0002b20e),
    .INIT_60(256'h022ffd2277f2b80e022ffd2070c20896022ffd2500022189022ffd206de01020),
    .INIT_61(256'h022ffd0bc022b80f022ffd206de20896022ffd2071622189022ffd2072001010),
    .INIT_62(256'h022ffd2074620896022ffd2075222202022ffd206dc2f01e022ffd206b601008),
    .INIT_63(256'h022ffd0bc3a2f01e022ffd206de01001022ffd2070c2b20f022ffd2071e2b40f),
    .INIT_64(256'h022ffd20714010a0022ffd250000b203022ffd206dc19801022ffd206b60982f),
    .INIT_65(256'h022ffd206e8208e4022ffd206e8208b7022ffd206de208d4022ffd2070601102),
    .INIT_66(256'h022ffd206b62fe0e022ffd0bc052fd0d022ffd206b62fc0c022ffd0bc0603f03),
    .INIT_67(256'h022ffd207e90be0e022ffd206dc0bd0d022ffd206b60bc0c022ffd0bc042ff0f),
    .INIT_68(256'h022ffd09502208d4022ffd206de01100022ffd206fe01020022ffd207220bf0f),
    .INIT_69(256'h022ffd227bf361aa022ffd207fb0d001022ffd3a7a80b001022ffd0d504208ee),
    .INIT_6A(256'h022ffd09f1f208c3022ffd09e1e208ab022ffd09d1d221ad022ffd09c1c22017),
    .INIT_6B(256'h022ffd10cb00b017022ffd14b061d000022ffd14b060b016022ffd0bb0220911),
    .INIT_6C(256'h022ffd2ff3b0b019022ffd13f001f000022ffd13e000b018022ffd13d001f000),
    .INIT_6D(256'h022ffd0bc3b0b01b022ffd2fc341f000022ffd2fd350b01a022ffd2fe361f000),
    .INIT_6E(256'h022ffd0bc350b01d022ffd206b61f000022ffd0bc360b01c022ffd206b61f000),
    .INIT_6F(256'h022ffd206dc1d002022ffd206b60b032022ffd0bc34361c9022ffd206b61f000),
    .INIT_70(256'h022ffd0d5042f03a022ffd206de11001022ffd206fe0b03a022ffd20700324cd),
    .INIT_71(256'h022ffd0bc343247a022ffd227dd1d001022ffd207fb0b032022ffd3a7c7208a5),
    .INIT_72(256'h022ffd01a04308fa022ffd0bf3b0d001022ffd0be360b001022ffd0bd3522008),
    .INIT_73(256'h022ffd09f072f034022ffd206280b016022ffd2067a321ff022ffd01b001d800),
    .INIT_74(256'h022ffd09d072f036022ffd206280b018022ffd09e072f035022ffd206280b017),
    .INIT_75(256'h022ffd00cd02f03c022ffd206b60b01a022ffd09c072f03b022ffd206280b019),
    .INIT_76(256'h022ffd00cf02f03e022ffd206b60b01c022ffd00ce02f03d022ffd206b60b01b),
    .INIT_77(256'h022ffd20712208ab022ffd20700208f1022ffd206dc2f03f022ffd206b60b01d),
    .INIT_78(256'h022ffd0d5040b134022ffd01c000b016022ffd206e820911022ffd206de208c3),
    .INIT_79(256'h022ffd206dc1e010022ffd206b60b135022ffd11c010b017022ffd14c001c010),
    .INIT_7A(256'h022ffd206de0b019022ffd207201e010022ffd207220b136022ffd250000b018),
    .INIT_7B(256'h022ffd206b60b13c022ffd09c0c0b01a022ffd2b03c1e010022ffd2b80c0b13b),
    .INIT_7C(256'h022ffd2b01c1e010022ffd206b60b13d022ffd09c0c0b01b022ffd2b02c1e010),
    .INIT_7D(256'h022ffd09c0c0b01d022ffd2b00c1e010022ffd206b60b13e022ffd09c0c0b01c),
    .INIT_7E(256'h022ffd2072a19801022ffd2500036211022ffd206dc1e010022ffd206b60b13f),
    .INIT_7F(256'h022ffd2072a20aad022ffd2072a221de022ffd2072a321ff022ffd2072a1d800),
    .INITP_00(256'h61a51039fc6e62cb9c200dfed57fe35bce36ed465530b584394da0b9af00ab01),
    .INITP_01(256'hb0128f908310a32685256ebf3b0c7ed14b7be11a2721ede8f1d62fbf25d65077),
    .INITP_02(256'h4acf7e68c94fcdffd7ea6a50ef66516a6ff8de69c4ffe6eaf87ce940455d2785),
    .INITP_03(256'h61f663f6ca707fcc4bfaface7b66f9ced74259fdecc6dd71447872e8e9e55a73),
    .INITP_04(256'h67c7d6dee1c0e0e2f8697df7c5c15ef465556df473dafa6ffe7159e77be9d876),
    .INITP_05(256'h7d4acb79c16ccad2e6524e644d7bf35e415b7e57e1caece0ce69794e68c065db),
    .INITP_06(256'h6e51655cea5fd3436be6ecc6d84350c64559527f6965f95de1f86acd6fca7355),
    .INITP_07(256'he7fbf860f8dd7c5d6652efc2e2dc7adcef45ef5bec50e04aef416a5cef5cef7e),
    .INITP_08(256'h6b6871606d7f65e765f5ed6df0616beff27bfcf4f0feea6ef279fc75f07f6bec),
    .INITP_09(256'hf1c869facb71efffdaea72fedde96a41f0786b7471e76b6565796a7ae174f0ff),
    .INITP_0A(256'hedf65bde74f3c44f6e56646ad350704c494d65fdf1d7d2f34dc1e042c3536c6d),
    .INITP_0B(256'h7bd5f4df4d6562d27369fa54cde9557c7045596a5465fffa7c594ec463fee95c),
    .INITP_0C(256'h4ceddbee537fd8e278fc7dca41e7ebcb62e25cd871fc724571f3cf5349d6faeb),
    .INITP_0D(256'he8c26ac667c665c67e71c14e79efc04bcf7863c7c976fcc553594968476cf4dd),
    .INITP_0E(256'h53567bcfc84c50cc524f5f6f7eecff6b5fe8ce4bf6754ad8f57fdbe571f4f9cf),
    .INITP_0F(256'h42cdd2dacd7965cdc95c4e4ac248ca43cb49ddec6a454a61654f51467b63f474),
