    localparam [35:0] init1FB = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init1FC = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init1FD = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init1FE = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init1FF = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init200 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init201 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init202 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init203 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init204 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init205 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init206 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init207 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init208 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init209 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init20A = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init20B = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init20C = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init20D = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init20E = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init20F = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init210 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init211 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init212 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init213 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init214 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init215 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init216 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init217 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init218 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init219 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init21A = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init21B = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init21C = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init21D = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init21E = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init21F = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init220 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init221 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init222 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init223 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init224 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init225 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init226 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init227 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init228 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init229 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init22A = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init22B = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init22C = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init22D = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init22E = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init22F = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init230 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init231 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init232 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init233 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init234 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init235 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init236 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init237 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init238 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init239 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init23A = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init23B = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init23C = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init23D = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init23E = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init23F = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init240 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init241 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init242 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init243 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init244 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init245 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init246 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init247 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init248 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init249 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init24A = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init24B = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init24C = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init24D = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init24E = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init24F = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init250 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init251 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init252 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init253 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init254 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init255 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init256 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init257 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init258 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init259 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init25A = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init25B = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init25C = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init25D = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init25E = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init25F = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init260 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init261 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init262 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init263 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init264 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init265 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init266 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init267 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init268 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init269 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init26A = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init26B = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init26C = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init26D = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init26E = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init26F = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init270 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init271 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init272 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init273 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init274 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init275 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init276 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init277 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init278 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init279 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init27A = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init27B = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init27C = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init27D = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init27E = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init27F = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init280 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init281 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init282 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init283 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init284 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init285 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init286 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init287 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init288 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init289 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init28A = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init28B = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init28C = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init28D = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init28E = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init28F = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init2F0 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init2F1 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init2F2 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init2F3 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init2F4 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init2F5 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init2F6 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init2F7 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init2F8 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init2F9 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init2FA = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init2FB = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init2FC = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init2FD = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init2FE = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init2FF = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init300 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init301 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init302 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init303 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init304 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init305 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init306 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init307 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init308 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init309 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init30A = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init30B = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init30C = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init30D = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init30E = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init30F = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init310 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init311 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init312 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init313 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init314 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init315 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init316 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init317 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init318 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init319 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init31A = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init31B = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init31C = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init31D = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init31E = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init31F = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init320 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init321 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init322 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init323 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init324 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init325 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init326 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init327 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init328 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init329 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init32A = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init32B = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init32C = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init32D = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init32E = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init32F = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init330 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init331 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init332 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init333 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init334 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init335 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init336 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init337 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init338 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init339 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init33A = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init33B = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init33C = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init33D = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init33E = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init33F = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init340 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init341 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init342 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init343 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init344 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init345 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init346 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init347 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init348 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init349 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init34A = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init34B = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init34C = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init34D = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init34E = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init34F = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init350 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init351 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init352 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init353 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init354 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init355 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init356 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init357 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init358 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init359 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init35A = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init35B = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init35C = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init35D = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init35E = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init35F = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init360 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init361 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init362 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init363 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init364 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init365 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init366 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init367 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init368 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init369 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init36A = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init36B = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init36C = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init36D = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init36E = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init36F = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init370 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init371 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init372 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init373 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init374 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init375 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init376 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init377 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init378 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init379 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init37A = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init37B = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init37C = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init37D = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init37E = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init37F = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init380 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init381 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init382 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init383 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init384 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init385 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init386 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
    localparam [35:0] init387 = {1'b1, 1'b1, 1'b1, 1'b1, 32'h00000000};
