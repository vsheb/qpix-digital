//defaulted to header of xcku040
`define x8_33554434
