    .INIT_00(256'h022ffc250001d000022ffc209280b016022ffc2b08e2f03a022ffc2bebb11001),
    .INIT_01(256'h022ffc208491f000022ffc208dc0b018022ffc01ccc1f000022ffc2079f0b017),
    .INIT_02(256'h022ffc2b10a1f000022ffc2b6490b01a022ffc207b21f000022ffc2079f0b019),
    .INIT_03(256'h022ffc2b6c91f000022ffc209280b01c022ffc2b08e1f000022ffc2bdfb0b01b),
    .INIT_04(256'h022ffc209282006d022ffc2b08e3602a022ffc2bebb1f000022ffc2b10a0b01d),
    .INIT_05(256'h022ffc208dc32193022ffc01cd81d002022ffc2079f0b002022ffc2500020076),
    .INIT_06(256'h022ffc208dc32193022ffc01ccc1d003022ffc2079f0b002022ffc208492007f),
    .INIT_07(256'h022ffc2b6490b032022ffc207b22085b022ffc2079f20700022ffc2084920088),
    .INIT_08(256'h022ffc20928325ba022ffc2b08e1d002022ffc2bdfb32542022ffc2b10a1d001),
    .INIT_09(256'h022ffc2b08e0bd10022ffc2bebb2f01e022ffc2b10a01001022ffc2b6c92200a),
    .INIT_0A(256'h022ffc01ce413e00022ffc2079f11d01022ffc250000bf12022ffc209280be11),
    .INIT_0B(256'h022ffc01cd803f03022ffc2079f2fe11022ffc208492fd10022ffc208dc13f00),
    .INIT_0C(256'h022ffc01ccc03007022ffc2079f0b00f022ffc2084920ba5022ffc208dc2ff12),
    .INIT_0D(256'h022ffc207b20be0e022ffc2079f030fc022ffc208490b03b022ffc208dc2f00f),
    .INIT_0E(256'h022ffc2b08e0b001022ffc2bdfb3626c022ffc2b10a1c0e0022ffc2b64903efc),
    .INIT_0F(256'h022ffc2bebb32248022ffc2b10a1d001022ffc2b6c932244022ffc209281d000),
    .INIT_10(256'h022ffc2b1c932250022ffc250001d003022ffc209283224c022ffc2b08e1d002),
    .INIT_11(256'h022ffc2092822253022ffc2b08e2093c022ffc2b47b207cd022ffc2b22a208e8),
    .INIT_12(256'h022ffc2b57b22253022ffc2b22a2093c022ffc2b489207d4022ffc25000208eb),
    .INIT_13(256'h022ffc2b5c922253022ffc250002093c022ffc20928207de022ffc2b08e208ee),
    .INIT_14(256'h022ffc209280b016022ffc2b08e2093c022ffc2b6bb207ea022ffc2b66a208f1),
    .INIT_15(256'h022ffc2b7bb0b018022ffc2b66a1f000022ffc2b6c90b017022ffc250001d000),
    .INIT_16(256'h022ffc2079f0b01a022ffc250001f000022ffc209280b019022ffc2b08e1f000),
    .INIT_17(256'h022ffc011010b01c022ffc010801f000022ffc2079f0b01b022ffc208551f000),
    .INIT_18(256'h022ffc2079f36265022ffc250001f000022ffc207c10b01d022ffc208b71f000),
    .INIT_19(256'h022ffc2079f2065e022ffc2084920713022ffc208dc206e1022ffc01c0e2226c),
    .INIT_1A(256'h022ffc01c1e2200a022ffc2079f206d2022ffc2500001004022ffc207a620724),
    .INIT_1B(256'h022ffc207a61d002022ffc2079f0b002022ffc2084920076022ffc208dc2006d),
    .INIT_1C(256'h022ffc2079f1d003022ffc208490b002022ffc208dc2007f022ffc01c0e32276),
    .INIT_1D(256'h022ffc01c2e2085b022ffc2079f20700022ffc2500020088022ffc207a632276),
    .INIT_1E(256'h022ffc207a62d010022ffc2079f01080022ffc208492b10f022ffc208dc2b80f),
    .INIT_1F(256'h022ffc2079f206d2022ffc2084901002022ffc208dc2d010022ffc01c1e01010),
    .INIT_20(256'h022ffc208492f032022ffc208dc01000022ffc01c0e2200a022ffc207a620713),
    .INIT_21(256'h022ffc0b00209017022ffc25000322b5022ffc207a60d004022ffc2079f0900e),
    .INIT_22(256'h022ffc3289009019022ffc1d0032f008022ffc3288e09018022ffc1d0022f007),
    .INIT_23(256'h022ffc228930901b022ffc208632f00a022ffc328920901a022ffc1d0042f009),
    .INIT_24(256'h022ffc0b0022b04e022ffc208762f033022ffc2289309016022ffc2086a2f00b),
    .INIT_25(256'h022ffc208dc09002022ffc01c0e3629b022ffc2079f1d00a022ffc250000300f),
    .INIT_26(256'h022ffc2079f1d00e022ffc2500022493022ffc2079f32492022ffc208490d002),
    .INIT_27(256'h022ffc2079f362a8022ffc208491d00b022ffc208dc22492022ffc01c1a3629e),
    .INIT_28(256'h022ffc2079f206a0022ffc208492dc01022ffc208dc03c0f022ffc01c0e0bc07),
    .INIT_29(256'h022ffc208dc22003022ffc01c262065e022ffc2079f20638022ffc2500020660),
    .INIT_2A(256'h022ffc208dc224b9022ffc01c1a206a6022ffc2079f362ac022ffc208491d00d),
    .INIT_2B(256'h022ffc208dc224a4022ffc01c0e20684022ffc2079f362b0022ffc208491d00f),
    .INIT_2C(256'h022ffc01019324bf022ffc250000d008022ffc2079f324bf022ffc208491d00c),
    .INIT_2D(256'h022ffc2b00a36492022ffc250000d020022ffc3e8b40900d022ffc1900122490),
    .INIT_2E(256'h022ffc2b00a09002022ffc2d108362bf022ffc2d0081d04f022ffc2b41909006),
    .INIT_2F(256'h022ffc250001d053022ffc2d10822493022ffc2d00832492022ffc2b2590d002),
    .INIT_30(256'h022ffc2dd080b202022ffc2dc082065e022ffc2b289206a2022ffc2b00a362cb),
    .INIT_31(256'h022ffc2b00a11301022ffc250002072b022ffc2df082071c022ffc2de0801300),
    .INIT_32(256'h022ffc09e081d052022ffc09d0822491022ffc09c08362c5022ffc2b2891c320),
    .INIT_33(256'h022ffc2d00909006022ffc2d10a206b5022ffc25000206a0022ffc09f08362e2),
    .INIT_34(256'h022ffc2df08206b5022ffc2de0820660022ffc2dd0836490022ffc2dc081d020),
    .INIT_35(256'h022ffc09c082066a022ffc2d00936490022ffc2d10a1d030022ffc2500009006),
    .INIT_36(256'h022ffc250003a490022ffc09f082062b022ffc09e0809006022ffc09d08206b5),
    .INIT_37(256'h022ffc2d009206b2022ffc2d10a20649022ffc0110200100022ffc010502d001),
    .INIT_38(256'h022ffc208c7362e6022ffc207c11d055022ffc2500022003022ffc2dc082065e),
    .INIT_39(256'h022ffc25000362ea022ffc207c71d044022ffc208c0224b9022ffc25000206a6),
    .INIT_3A(256'h022ffc2089536311022ffc250001d04e022ffc208f4224a4022ffc2079f20684),
    .INIT_3B(256'h022ffc208f41d020022ffc2089b09006022ffc25000206b5022ffc208f420698),
    .INIT_3C(256'h022ffc250002064e022ffc208f40120a022ffc208a520660022ffc2500036490),
    .INIT_3D(256'h022ffc0bf0f2fc0a022ffc208b72fb09022ffc011002fa08022ffc010203a490),
    .INIT_3E(256'h022ffc208e52064e022ffc0bc0c01201022ffc0bd0d2fe33022ffc0be0e2fd0b),
    .INIT_3F(256'h022ffc0110114a06022ffc0108014a06022ffc208e814a06022ffc250003a490),
    .INIT_40(256'h022ffc208d50bd0a022ffc011000bc09022ffc010000bb08022ffc208b714a06),
    .INIT_41(256'h022ffc208eb20624022ffc2500020624022ffc207f80bf33022ffc208e50be0b),
    .INIT_42(256'h022ffc208b72fb08022ffc011012fa07022ffc0108020624022ffc2089520624),
    .INIT_43(256'h022ffc208e52ff33022ffc208d52fe0b022ffc011002fd0a022ffc010042fc09),
    .INIT_44(256'h022ffc2089b206a4022ffc208ee3637e022ffc250001d054022ffc20804224d0),
    .INIT_45(256'h022ffc0100836490022ffc208b71d020022ffc0110109006022ffc01080206b5),
    .INIT_46(256'h022ffc208153a490022ffc208e52064e022ffc208d50120a022ffc0110020660),
    .INIT_47(256'h022ffc010802fd0b022ffc208a52fc0a022ffc208f12fb09022ffc250002fa08),
    .INIT_48(256'h022ffc011003a490022ffc0100c2064e022ffc208b701201022ffc011012fe33),
    .INIT_49(256'h022ffc2500014a06022ffc2082a14a06022ffc208e514a06022ffc208d53a490),
    .INIT_4A(256'h022ffc250000bb08022ffc369280ba07022ffc0d0082fa07022ffc0900e14a06),
    .INIT_4B(256'h022ffc250000bf33022ffc3292c0be0b022ffc0d0020bd0a022ffc0900e0bc09),
    .INIT_4C(256'h022ffc2500020624022ffc3293020624022ffc0d00220624022ffc0900f20624),
    .INIT_4D(256'h022ffc250002fd0a022ffc329342fc09022ffc0d0022fb08022ffc090102fa07),
    .INIT_4E(256'h022ffc250002fb3f022ffc329382fa3e022ffc0d0022ff33022ffc090112fe0b),
    .INIT_4F(256'h022ffc2f11732341022ffc2f1160df08022ffc0110032360022ffc370011df0c),
    .INIT_50(256'h022ffc2f11b2061d022ffc2f11a2fa13022ffc2f1190ba33022ffc2f11822490),
    .INIT_51(256'h022ffc2b6c92fc0c022ffc010a22061d022ffc2f11d2061d022ffc2f11c2061d),
    .INIT_52(256'h022ffc2095220aa0022ffc110012ff0f022ffc2b00b2fe0e022ffc2b00a2fd0d),
    .INIT_53(256'h022ffc3694a0bf12022ffc1d0ff0be11022ffc209b10bd10022ffc209572065e),
    .INIT_54(256'h022ffc09d0820638022ffc09c0800cf0022ffc250002066a022ffc3700020682),
    .INIT_55(256'h022ffc1d0d020638022ffc2500000cd0022ffc09f0820638022ffc09e0800ce0),
    .INIT_56(256'h022ffc001f020649022ffc329822063f022ffc1d0d12063f022ffc3296d0bc3f),
    .INIT_57(256'h022ffc001d022490022ffc209a020638022ffc001e00bc3e022ffc209a0206b2),
    .INIT_58(256'h022ffc011002061d022ffc209a02fe13022ffc001c02061d022ffc209a02061d),
    .INIT_59(256'h022ffc2f12e2fd11022ffc2f12c2fc10022ffc2f12a03e03022ffc2f1282061d),
    .INIT_5A(256'h022ffc2f12f0bf0c022ffc2f12d2065e022ffc2f12b20ba5022ffc2f1292fe12),
    .INIT_5B(256'h022ffc001e020638022ffc209a00bc0f022ffc001f00bd0e022ffc250000be0d),
    .INIT_5C(256'h022ffc001c020638022ffc209a000ce0022ffc001d020638022ffc209a000cd0),
    .INIT_5D(256'h022ffc2f52c2063f022ffc2f62a0bc3f022ffc2f72820638022ffc209a000cf0),
    .INIT_5E(256'h022ffc016000bc3e022ffc01500206b2022ffc0140020649022ffc2f42e2063f),
    .INIT_5F(256'h022ffc2f52d3639c022ffc2f62b1d058022ffc2f72922490022ffc0170020638),
    .INIT_60(256'h022ffc209a0206ac022ffc001f03e39c022ffc2296c0d004022ffc2f42f09002),
    .INIT_61(256'h022ffc209a036490022ffc001d01d020022ffc209a009006022ffc001e0206b5),
    .INIT_62(256'h022ffc0310f3a490022ffc001702064e022ffc209a001208022ffc001c020660),
    .INIT_63(256'h022ffc0310f2fc36022ffc001602fb35022ffc037f02fa34022ffc2f1292065e),
    .INIT_64(256'h022ffc0310f0be36022ffc001500bd35022ffc036f00bc34022ffc2f12b2fd3b),
    .INIT_65(256'h022ffc0310f205f5022ffc0014001b00022ffc035f001a01022ffc2f12d0bf3b),
    .INIT_66(256'h022ffc2f12822490022ffc0110020638022ffc034f009c07022ffc2f12f205ed),
    .INIT_67(256'h022ffc2296c206b5022ffc2f12e2069e022ffc2f12c3640f022ffc2f12a1d051),
    .INIT_68(256'h022ffc1450020660022ffc1410036490022ffc144001d020022ffc1410009006),
    .INIT_69(256'h022ffc147002fa08022ffc141003a490022ffc146002064e022ffc141000120a),
    .INIT_6A(256'h022ffc145002fe33022ffc141002fd0b022ffc144002fc0a022ffc141002fb09),
    .INIT_6B(256'h022ffc1470014a06022ffc141003a490022ffc146002064e022ffc1410001201),
    .INIT_6C(256'h022ffc0b9290bb08022ffc0b82814a06022ffc0017014a06022ffc2500014a06),
    .INIT_6D(256'h022ffc01b000bf33022ffc20a7c0be0b022ffc20a5e0bd0a022ffc20a520bc09),
    .INIT_6E(256'h022ffc0ba2620624022ffc14b0020624022ffc14a0e20624022ffc0ba2520624),
    .INIT_6F(256'h022ffc14b002fd0a022ffc14a002fc09022ffc14b002fb08022ffc14a002fa07),
    .INIT_70(256'h022ffc062b0323d1022ffc0b2171df0c022ffc14b002ff33022ffc14a002fe0b),
    .INIT_71(256'h022ffc14a002ff13022ffc14b0022490022ffc14a00323c7022ffc2f2170df08),
    .INIT_72(256'h022ffc14a002061d022ffc14b002061d022ffc14a002061d022ffc14b002061d),
    .INIT_73(256'h022ffc0ba272ff0f022ffc14b002fe0e022ffc14a002fd0d022ffc14b002fc0c),
    .INIT_74(256'h022ffc14b002fe13022ffc14a002061d022ffc14b002061d022ffc14a00223e6),
    .INIT_75(256'h022ffc06b202fc10022ffc0b21603e03022ffc14b002061d022ffc14a002061d),
    .INIT_76(256'h022ffc0b92b0b105022ffc0b82a0b004022ffc001602fe12022ffc2fb162fd11),
    .INIT_77(256'h022ffc01b001ae20022ffc20a7c1ad10022ffc20a5e18c00022ffc20a520b206),
    .INIT_78(256'h022ffc0ba2603407022ffc14b000b40f022ffc14a0e20ba5022ffc0ba253e490),
    .INIT_79(256'h022ffc14b000b013022ffc14a0020887022ffc14b00223e6022ffc14a002f40f),
    .INIT_7A(256'h022ffc062b0323f3022ffc0b2191d001022ffc14b00323f0022ffc14a001d000),
    .INIT_7B(256'h022ffc14a00323f9022ffc14b001d003022ffc14a00323f6022ffc2f2191d002),
    .INIT_7C(256'h022ffc14a00208eb022ffc14b00223fb022ffc14a00207cd022ffc14b00208e8),
    .INIT_7D(256'h022ffc0ba27207de022ffc14b00208ee022ffc14a00223fb022ffc14b00207d4),
    .INIT_7E(256'h022ffc14b002065e022ffc14a00207ea022ffc14b00208f1022ffc14a00223fb),
    .INIT_7F(256'h022ffc06b2009f0802d0030b2180125d0010ff14b002b6c902bff014a002b00a),
    .INITP_00(256'h4a455fc67cd355c27cd255c8494971c5ecc1515dccc7d6ddccfac6d951435160),
    .INITP_01(256'hf75ceb58504940cc40c04cf0d157dc66c8c9d76ad550d1d3497dcbfc40c7df5c),
    .INITP_02(256'hf4e558d3db42c45178d0675143ced5c773dd4c48cbcb6c5e53ce784e46574bc7),
    .INITP_03(256'hd9cdedcd4f5a53f5d25f48d547cbf8dfc25546f4d0d94055d44e78c2c8427e54),
    .INITP_04(256'h4dde6bc3455cd94ce244c35244c9e4d2e6d6d4f649e84e75c642d7c7cb724ed6),
    .INITP_05(256'hd5c87e75fbc06a47f0cd46c45d40515e6b54c358e0d9cbdd625a56c354c3f842),
    .INITP_06(256'he5c2e46959ffc55af0755dd0fbd34f6f7dc744e2434b6f60fdc474d5dc70eb77),
    .INITP_07(256'h76ed6359ff4eeaeb5cc37d434d7cd0d8ed58c876c95ee958d36eff4764e3d670),
    .INITP_08(256'h764ce55b69ff79e540cdec6f4af355e569e1744040e0e9dce64eeb63627c505c),
    .INITP_09(256'hefe562d4d5cf4679524ccb6d4e47d361d8c7cc6f55fc477f4afbf86a7fc95dea),
    .INITP_0A(256'h4670447ece77ecf776447052d47f4148d7f5e8ed75ed607ff2ea6d77eaeae2f8),
    .INITP_0B(256'hd5d4e2e15d4bed64dc40e4f8c4715a72db6fd4d2e2e1f0e67e6b7beaef6a4bff),
    .INITP_0C(256'hd4e765e8796047f04e74f3fa5e6bf570536854fdd7ecf941eec7e655f3c3ddee),
    .INITP_0D(256'hd3fbd77ed3cff6527c7c78f24f69eb4ac85aec48f0d25ad6d95aec49e5dbded3),
    .INITP_0E(256'h7a73606549fee0e0c9f9486bdd6b487fde5670dd6b486b48f3db6078eced5a70),
    .INITP_0F(256'h54f881714562d4f4c2daf446fcd768d967d6e0ebe3e8c0f3cefc5c694749ead1),
