    .INIT_00(256'h00000014a001fb0100000014b001dac000000014a003241b00000014b001fb01),
    .INIT_01(256'h0000000ba273241b00000014b001fb0200000014a001da0000000014b003241b),
    .INIT_02(256'h00000014b001da8000000014a003241b00000014b001fb0200000014a001da20),
    .INIT_03(256'h00000006b201fb020000000b2181daa000000014b003241b00000014a001fb02),
    .INIT_04(256'h0000000b92d3241b0000000b82c1fb02000000001501dac00000002fb183241b),
    .INIT_05(256'h00000001b001dae000000020a8c3241b00000020a6e1fb0300000020a621da00),
    .INIT_06(256'h0000000ba262071600000014b002242d00000014a0e3241b0000000ba251fb03),
    .INIT_07(256'h00000014b002090f00000014a00001b000000014b00000a000000014a00208d1),
    .INIT_08(256'h000000062b000cf00000000b21b00bc000000014b002091f00000014a00208f2),
    .INIT_09(256'h00000014a0000cd000000014b00206f000000014a0000ce00000002f21b206f0),
    .INIT_0A(256'h00000014a00208e000000014b00206f000000014a0000cb000000014b00206f0),
    .INIT_0B(256'h0000000ba272200800000014b00207b500000014a002071600000014b002242d),
    .INIT_0C(256'h00000014b002012800000014a00208d100000014b002071600000014a0020752),
    .INIT_0D(256'h00000006b202b80f0000000b21a2b40f00000014b002b20f00000014a00208e0),
    .INIT_0E(256'h0000000b92f220080000000b82e207b500000000140207870000002fb1a01002),
    .INIT_0F(256'h00000001b00208e000000020a8c2012800000020a6e208d100000020a6220716),
    .INIT_10(256'h0000000ba260100000000014b002b80f00000014a0e2b40f0000000ba252b20f),
    .INIT_11(256'h00000014b00207a300000014a002f03200000014b000100100000014a002f01e),
    .INIT_12(256'h000000062b0224bf0000000b21d2071800000014b002071c00000014a002073c),
    .INIT_13(256'h00000014a002b40f00000014b002b20f00000014a00208d10000002f21d20716),
    .INIT_14(256'h00000014a00207a300000014b002f03200000014a000100200000014b002b80f),
    .INIT_15(256'h0000000ba270bc3300000014b002071800000014a002075000000014b0022500),
    .INIT_16(256'h00000014b002076a00000014a002070100000014b00206f700000014a00206f7),
    .INIT_17(256'h00000006b20206f00000000b21c0bc0a00000014b00206f000000014a000bc0b),
    .INIT_18(256'h00000001b00206f000000001a000bc0800000025000206f00000002fb1c0bc09),
    .INIT_19(256'h00000014a00090020000000d8ff2071600000014a00206f00000000d1ff0bc07),
    .INIT_1A(256'h00000014b00010100000000daff208d100000014a003246e0000000d9ff0d008),
    .INIT_1B(256'h00000001a0020787000000002000100000000025000220080000002fb2520787),
    .INIT_1C(256'h00000014a040bb0800000014a040ba0700000014a00220080000000d1ff207b5),
    .INIT_1D(256'h00000014a040bf3300000014a040be0b00000014a040bd0a00000014a040bc09),
    .INIT_1E(256'h00000020a7f3247f000000022a01d00c00000014a040300f00000014a04000f0),
    .INIT_1F(256'h00000000a80000a000000025000224ba0000002f2263247f000000062b00d008),
    .INIT_20(256'h00000014a06206d500000014b00206d500000014a062f01400000000b900301f),
    .INIT_21(256'h00000014a061d05d00000014b000307f00000014a06000b000000014b00206d5),
    .INIT_22(256'h000000250000300f00000014b000b03300000014a062f01500000014b003e4ba),
    .INIT_23(256'h00000001b003249900000001a000d0080000000038032490000000002101d00c),
    .INIT_24(256'h00000014a002f0130000000d2ff03003000000033011400e000000032aa000e0),
    .INIT_25(256'h00000014b08206d50000000daff364ba00000014a001c0100000000d3ff0b102),
    .INIT_26(256'h000000032cc2f01300000001a0003003000000003800b03300000000210364a8),
    .INIT_27(256'h0000000d3ff206d500000014a00364ba0000000d2ff1c010000000033020b102),
    .INIT_28(256'h000000002102ff0f00000014b082fe0e0000000daff2fd0d00000014a002fc0c),
    .INIT_29(256'h00000003304224b7000000032f0324ba00000001a001df010000000038003f07),
    .INIT_2A(256'h00000014a002fe120000000d3ff2fd1100000014a002fc100000000d2ff03e03),
    .INIT_2B(256'h0000002500018c000000002fb270b20600000014b080b1050000000daff0b004),
    .INIT_2C(256'h0000000110020bec0000000100c3e4ba000000008401ae20000000009501ad10),
    .INIT_2D(256'h0000001900120935000000131002f40f00000014808034070000001490e0b40f),
    .INIT_2E(256'h000000019ff0100000000036abe208e00000001d1002093900000036ab4206ba),
    .INIT_2F(256'h00000036ac40900f0000000d5082200800000025000207b5000000018ff20787),
    .INIT_30(256'h000000250003617c000000018ff0d020000000019ff3617c000000011020d040),
    .INIT_31(256'h000000000400d080000000001500900e0000003ead1361770000001d1030d080),
    .INIT_32(256'h000000140080d0200000001410e36170000000118010d040000000018ff36173),
    .INIT_33(256'h000000011040900e0000000190b3616a000000118080d0100000003eac93616d),
    .INIT_34(256'h000000198182f033000000008400901600000000950324d9000000250000d004),
    .INIT_35(256'h000000019ff324e8000000011021d00e0000003eada0300f0000001b9052b04e),
    .INIT_36(256'h0000000381f364bf000000001800d020000000250000900d000000018ff224bf),
    .INIT_37(256'h000000149001d05300000014106324e8000000149001d0490000001410609006),
    .INIT_38(256'h00000000080207be0000000110220716000000149002075a00000014106364bf),
    .INIT_39(256'h00000014006224bf0000001400620718000000140062071c00000000a902073c),
    .INIT_3A(256'h00000014a002011e00000014006208d100000014a00207160000001400620746),
    .INIT_3B(256'h00000036af22d0030000001d90b2f0320000003d000010000000001da5d208e0),
    .INIT_3C(256'h000000250002200800000001104207b50000003aaf4207870000001d81401000),
    .INIT_3D(256'h000000370010106000000025000208e00000003aaf22011e0000001d808208d1),
    .INIT_3E(256'h0000000b40e2d0030000000b30d2f0320000000b20c0100000000020bd12077b),
    .INIT_3F(256'h0000001450e2200800000003403207b500000000540207870000000ba0f01000),
    .INIT_40(256'h000000007a02fd100000000360701f00000000006a001e000000001450e01d00),
    .INIT_41(256'h0000001470e2fd1e0000001470e01d010000001470e2ff120000001470e2fe11),
    .INIT_42(256'h000000008203251200000001e001d0ff00000001d000b00f0000000370320bec),
    .INIT_43(256'h00000032b5b209350000001d6032f00f00000032b33030070000001d6020b00f),
    .INIT_44(256'h00000001a000d004000000019000900e00000032b912219e0000001d6042094c),
    .INIT_45(256'h00000032b1f2b04e0000001ce402f03300000036b18090160000001cd303251b),
    .INIT_46(256'h00000013a000b004000000139003252d000000108f01d00e00000009f080300f),
    .INIT_47(256'h00000001d000be1100000022b140bd1000000013e000b20600000011d010b105),
    .INIT_48(256'h00000032b291ee100000001cd501cd000000000bf3103f010000000be300bf12),
    .INIT_49(256'h00000011d0113e0000000013a0011d01000000129f03252d000000108e01ef20),
    .INIT_4A(256'h00000003a032ff120000002f9112fe110000002f8102fd1000000022b2213f00),
    .INIT_4B(256'h00000004a00208e0000000140062011e00000014006208d10000000b00222506),
    .INIT_4C(256'h0000000bd30207870000002500001000000000370002d1030000002fa1201000),
    .INIT_4D(256'h00000001a001d001000000019000b01e0000000b237220080000000be31207b5),
    .INIT_4E(256'h000000108d00b51700000032b400b4160000001cf200120000000001f0036590),
    .INIT_4F(256'h00000022b390421000000011f012f91700000013a002f816000000129e020ab0),
    .INIT_50(256'h00000032b492f8180000001cf5020ab00000000b23c0b51900000001f000b418),
    .INIT_51(256'h00000011f010b51b00000013a000b41a0000001390004210000000108202f919),
    .INIT_52(256'h00000032b51042100000001cf302f91b00000001f002f81a00000022b4220ab0),
    .INIT_53(256'h00000011f012f81c0000001380020ab0000000139000b51d000000118020b41c),
    .INIT_54(256'h00000003a03325610000002f9110d2020000002f8100421000000022b4a2f91d),
    .INIT_55(256'h00000004a002083e0000001400620853000000140062f21e0000000b00201202),
    .INIT_56(256'h0000000bd30324f4000000250001d001000000370000b0320000002fa122084b),
    .INIT_57(256'h000000019000502000000001800207750000000b237325120000000be311d002),
    .INIT_58(256'h00000032b6920cc80000001cf202f21e00000001f000120400000001a00225d1),
    .INIT_59(256'h00000011f012f11500000013a002f014000000129e00b117000000108d00b016),
    .INIT_5A(256'h0000001df000b01800000003ff0346ba0000000bf391f1ff00000022b621d0ff),
    .INIT_5B(256'h0000001df021d0ff0000000b23c2f11500000001f002f01400000032b760b119),
    .INIT_5C(256'h00000013a000b11b000000139000b01a00000010820346ba00000032b761f1ff),
    .INIT_5D(256'h0000000b2381f1ff00000001f001d0ff00000022b6f2f11500000011f012f014),
    .INIT_5E(256'h000000139002f014000000108200b11d00000032b7f0b01c0000001cf50346ba),
    .INIT_5F(256'h00000001f00346ba00000022b781f1ff00000011f011d0ff00000013a002f115),
    .INIT_60(256'h0000001390020939000000118013658400000032b871d0000000001cf300b032),
    .INIT_61(256'h0000002f8102084b00000022b802087b00000011f012083e0000001380020853),
    .INIT_62(256'h000000140061d0020000000b002324f400000003a031d0010000002f9110b032),
    .INIT_63(256'h00000037000225d10000002fa12030df00000004a00207750000001400632512),
    .INIT_64(256'h0000000b237207580000000be312073a0000000bd303659d000000250001d008),
    .INIT_65(256'h00000001f000b03200000001a00208230000000190020716000000018002073a),
    .INIT_66(256'h000000129e005020000000108d02077500000032b9f324f40000001cf201d001),
    .INIT_67(256'h0000000bf392073600000022b98365aa00000011f011d01000000013a00225d1),
    .INIT_68(256'h00000001f002082300000032bac207160000001df002076400000003ff02075e),
    .INIT_69(256'h000000108202077500000032bac324f40000001df021d0010000000b23c0b032),
    .INIT_6A(256'h00000022ba5365b700000011f011d02000000013a00225d10000001390005020),
    .INIT_6B(256'h0000001cf00207160000000b037207640000000b2382075e00000001f0020736),
    .INIT_6C(256'h00000013a00324f4000000139001d001000000108200b03200000032bb620823),
    .INIT_6D(256'h0000000b2031d04000000001f00225d100000022bae030df00000011f0120775),
    .INIT_6E(256'h0000001390020764000000108202075e00000032bbf207360000001cf50365c4),
    .INIT_6F(256'h00000001f001d00100000022bb80b03200000011f012082300000013a0020716),
    .INIT_70(256'h00000013900225d100000011801030df00000032bc7207750000001cf30324f4),
    .INIT_71(256'h0000002f8102075200000022bc02075800000011f0136017000000138001d080),
    .INIT_72(256'h000000140060b0320000000b0022082300000003a03207160000002f9112074e),
    .INIT_73(256'h00000037000030df0000002fa122077500000004a00324f4000000140061d001),
    .INIT_74(256'h0000002f50320787000000095080100800000020be52077b00000025000225d1),
    .INIT_75(256'h0000002f6053663f0000002f5041d004000000096080b01e0000000950822008),
    .INIT_76(256'h0000002f631206830000002f5303262a000000096080d0040000000950809002),
    .INIT_77(256'h0000002f638011b30000002f53701e400000000960801f0a00000009508206a9),
    .INIT_78(256'h0000002f6062df0a0000002f53c09d070000000960820663000000095080120b),
    .INIT_79(256'h00000001100365eb000000016071ce10000000015ef2dd08000000250002de09),
    .INIT_7A(256'h0000002500011e010000002d10b225ee0000002d60a365eb0000002d5091cf20),
    .INIT_7B(256'h0000000b9110b1170000000b8100b01600000020bd1225e10000003700113f00),
    .INIT_7C(256'h0000002fa361f1ff0000002f9351d0ff0000002f8342f1150000000ba122f014),
    .INIT_7D(256'h0000000b4310d0ff0000000b330012000000000bd372066b00000001200325fa),
    .INIT_7E(256'h0000003ac030b1190000001ba000b0180000001a9402f2200000001883014200),
    .INIT_7F(256'h0000002fa361f1ff0000002f9351d0ff0000002f8342f115000000112012f014),
    .INITP_00(256'haf82258baea08f3c91188811319c01173e1eb60135952210b0229ab6073e9524),
    .INITP_01(256'h0d9a811abc97950e2a12a90b348bb21ca6b291a00bb191b110b113949c162607),
    .INITP_02(256'had96b18b3b983112aab699251b3217360ba98b10051130993811321aad361134),
    .INITP_03(256'h26a48e121c351a98909919121d9783943236218f382f98370291920f94a83090),
    .INITP_04(256'hbc849c0f31a2b4b2a3201ebd1805141d9a313dbea4b29cb2022d083e9a3e1f12),
    .INITP_05(256'h9bbc3314b2b6a0a03118b7010db70db0bf9a22b68b2f00159039be39373d2208),
    .INITP_06(256'h06310da236182700371e3381918aad371bb62da286b828063e9faa32209aa207),
    .INITP_07(256'h1d3ab03598289218a8a9893f21090e391f07b122178e911606901627328e9ca7),
    .INITP_08(256'h09a99aaa34390e921c3ca991b0212013a01f8f06250694a53338bcb7129cbe1f),
    .INITP_09(256'h3090aa9d0fbeafa2a3bb1e8893302e35a0128ebb8a2c952bb1321c820b332586),
    .INITP_0A(256'h2e9781999b24b3abaa8711a71e398b029c053ca2b82e2e980c36b29420949ab6),
    .INITP_0B(256'hba8094303980328a85258d0a373e0b311697bbbd9190bf0684be8a0ebe2739ae),
    .INITP_0C(256'hbc841ead9606adb531af331b038307a02aafbd1985a18ab3948893002dbeb4bf),
    .INITP_0D(256'ha58918b7bd0fb6960ea88a84392780a0bd250038151dad2d84ad9693a9239794),
    .INITP_0E(256'habb39c82a6bc0414a4b98895b0838529a9b1b48317349db584b89d0b2a3806b2),
    .INITP_0F(256'hbca48d2a13169eaa8bbf8f15bca48d3a34838231b5b887090cb52db23d32008b),
