    .INIT_00(256'h0000000b92d206380000000b82c09c080000000015009d080000002fb1809e08),
    .INIT_01(256'h00000001b002063800000020a7c00ce000000020a5e2063800000020a5200cd0),
    .INIT_02(256'h0000000ba261920100000014b002065e00000014a0e206380000000ba2500cf0),
    .INIT_03(256'h00000014b001d05000000014a002249100000014b002085b00000014a00363ff),
    .INIT_04(256'h000000062b0090060000000b21b206b500000014b002069c00000014a0036492),
    .INIT_05(256'h00000014a000120200000014b002066000000014a00364900000002f21b1d020),
    .INIT_06(256'h00000014a002061d00000014b002061d00000014a003a49000000014b002064e),
    .INIT_07(256'h0000000ba272061d00000014b002061d00000014a002fb1300000014b002061d),
    .INIT_08(256'h00000014b0003b0300000014a003645800000014b000d04000000014a0009002),
    .INIT_09(256'h00000006b201da200000000b21a3245800000014b001fb0000000014a001da00),
    .INIT_0A(256'h0000000b92f1fb000000000b82e1da8000000000140324580000002fb1a1fb00),
    .INIT_0B(256'h00000001b003245800000020a7c1fb0000000020a5e1daa000000020a5232458),
    .INIT_0C(256'h0000000ba261dae000000014b003245800000014a0e1fb000000000ba251dac0),
    .INIT_0D(256'h00000014b001fb0100000014a001da2000000014b003245800000014a001fb00),
    .INIT_0E(256'h000000062b0324580000000b21d1fb0100000014b001da8000000014a0032458),
    .INIT_0F(256'h00000014a001dac000000014b003245800000014a001fb010000002f21d1daa0),
    .INIT_10(256'h00000014a001fb0200000014b001da0000000014a003245800000014b001fb01),
    .INIT_11(256'h0000000ba273245800000014b001fb0200000014a001da2000000014b0032458),
    .INIT_12(256'h00000014b001daa000000014a003245800000014b001fb0200000014a001da80),
    .INIT_13(256'h00000006b201fb020000000b21c1dac000000014b003245800000014a001fb02),
    .INIT_14(256'h00000001b003245800000001a001fb03000000250001da000000002fb1c32458),
    .INIT_15(256'h00000014a00224900000000d8ff3245800000014a001fb030000000d1ff1dae0),
    .INIT_16(256'h00000014b001d0000000000daff0b01300000014a00208870000000d9ff2065e),
    .INIT_17(256'h00000001a001d0020000000020032468000000250001d0010000002fb2532463),
    .INIT_18(256'h00000014a04000a000000014a043247a00000014a001d0030000000d1ff32470),
    .INIT_19(256'h00000014a042248500000014a04208e200000014a04208b700000014a04001b0),
    .INIT_1A(256'h00000020a6f000a0000000022a02079f00000014a042085500000014a042079f),
    .INIT_1B(256'h00000000a802248500000025000208e20000002f226208b7000000062b0001b0),
    .INIT_1C(256'h00000014a062085500000014b002079f00000014a062085500000000b902079f),
    .INIT_1D(256'h00000014a06208b700000014b00001b000000014a06000a000000014b002079f),
    .INIT_1E(256'h000000250002085500000014b002079f00000014a062248500000014b00208e2),
    .INIT_1F(256'h00000001b002085500000001a002079f0000000038020855000000002102079f),
    .INIT_20(256'h00000014a00208b70000000d2ff001b000000003301000a0000000032aa2079f),
    .INIT_21(256'h00000014b08206380000000daff00cf000000014a0000bc00000000d3ff208e2),
    .INIT_22(256'h000000032cc2063800000001a0000cd000000000380206380000000021000ce0),
    .INIT_23(256'h0000000d3ff2249000000014a002085b0000000d2ff206380000000330200cb0),
    .INIT_24(256'h000000002102069a00000014b082200a0000000daff2071300000014a002065e),
    .INIT_25(256'h000000033040b002000000032f02007600000001a002006d000000003802065e),
    .INIT_26(256'h00000014a000b0020000000d3ff2007f00000014a003249f0000000d2ff1d002),
    .INIT_27(256'h000000250002085b0000002fb272008800000014b083249f0000000daff1d003),
    .INIT_28(256'h0000000b30d2200a0000000b20c2071300000020b7a206d20000003700101002),
    .INIT_29(256'h000000034030b00200000000540200760000000ba0f2006d0000000b40e2065e),
    .INIT_2A(256'h000000036070b002000000006a02007f0000001450e324af0000001450e1d002),
    .INIT_2B(256'h0000001470e2085b0000001470e200880000001470e324af000000007a01d003),
    .INIT_2C(256'h00000001e002f03200000001d0001001000000037032f01e0000001470e01000),
    .INIT_2D(256'h0000001d6032066000000032adc206640000001d6022068400000000820206ee),
    .INIT_2E(256'h000000019000100200000032b3a208870000001d6042065e00000032b0422542),
    .INIT_2F(256'h0000001ce402069800000036ac12258f0000001cd30206ee00000001a002f032),
    .INIT_30(256'h000000139002063f000000108f02063f00000009f080bc3300000032ac820660),
    .INIT_31(256'h00000022abd2063800000013e000bc0b00000011d01206b200000013a0020649),
    .INIT_32(256'h0000001cd50206380000000bf310bc090000000be302063800000001d000bc0a),
    .INIT_33(256'h00000013a0020638000000129f00bc07000000108e02063800000032ad20bc08),
    .INIT_34(256'h0000002f911324d80000002f8100d00800000022acb0900200000011d012065e),
    .INIT_35(256'h000000140062200a00000014006206d20000000b0130101000000003a0320887),
    .INIT_36(256'h000000250002200a00000037000207130000002fa12206d200000004a0001000),
    .INIT_37(256'h000000019000bd0a0000000b2370bc090000000be310bb080000000bd300ba07),
    .INIT_38(256'h00000032ae90300f0000001cf20000f000000001f000bf3300000001a000be0b),
    .INIT_39(256'h00000011f01324e900000013a000d008000000129e0324e9000000108d01d00c),
    .INIT_3A(256'h0000001cf502f0140000000b23c0301f00000001f00000a000000022ae22253d),
    .INIT_3B(256'h00000013a00000b0000000139002061d000000108202061d00000032af22061d),
    .INIT_3C(256'h0000001cf302f01500000001f003e53d00000022aeb1d05d00000011f010307f),
    .INIT_3D(256'h00000013800324fa000000139001d00c000000118020300f00000032afa0b033),
    .INIT_3E(256'h0000002f9111400e0000002f810000e000000022af33250300000011f010d008),
    .INIT_3F(256'h000000140061c010000000140060b1130000000b0132f01300000003a0303003),
    .INIT_40(256'h000000250000b03300000037000365120000002fa122061d00000004a003653d),
    .INIT_41(256'h000000018001c0100000000b2370b1130000000be312f0130000000bd3003003),
    .INIT_42(256'h0000001cf202fd0d00000001f002fc0c00000001a002061d000000019003653d),
    .INIT_43(256'h00000013a001df01000000129e003f07000000108d02ff0f00000032b122fe0e),
    .INIT_44(256'h00000003ff02fc100000000bf3903e0300000022b0b2252100000011f013253d),
    .INIT_45(256'h0000000b23c0b10500000001f000b00400000032b1f2fe120000001df002fd11),
    .INIT_46(256'h000000139001ae20000000108201ad1000000032b1f18c000000001df020b206),
    .INIT_47(256'h00000001f000340700000022b180b40f00000011f0120ba500000013a003e53d),
    .INIT_48(256'h000000108203252a00000032b281d0000000001cf500b0130000000b2382f40f),
    .INIT_49(256'h00000022b213253400000011f011d00200000013a003252f000000139001d001),
    .INIT_4A(256'h00000011801207cd00000032b30208e80000001cf303253900000001f001d003),
    .INIT_4B(256'h00000022b29208eb00000011f012253d00000013800208fd0000001390020602),
    .INIT_4C(256'h0000000b0132253d00000003a03209070000002f911206020000002f810207d4),
    .INIT_4D(256'h0000002fa122091200000004a002060200000014006207de00000014006208ee),
    .INIT_4E(256'h0000000be31206020000000bd30207ea00000025000208f1000000370002253d),
    .INIT_4F(256'h00000001a00206d20000000190001000000000018002085b0000000b2372091d),
    .INIT_50(256'h000000108d00d00800000032b48090110000001cf202200a00000001f0020713),
    .INIT_51(256'h00000022b413610700000011f010d08000000013a000900e000000129e036097),
    .INIT_52(256'h00000032b55360ff0000001df000d02000000003ff0361030000000bf390d040),
    .INIT_53(256'h00000032b550d0040000001df020900e0000000b23c360fb00000001f000d010),
    .INIT_54(256'h00000011f012b04e00000013a002f03300000013900090160000001082032558),
    .INIT_55(256'h0000000b037225420000000b2383256c00000001f001d00e00000022b4e0300f),
    .INIT_56(256'h0000001390009006000000108203654200000032b5f0d0200000001cf000900d),
    .INIT_57(256'h00000001f003654200000022b571d05300000011f013256c00000013a001d049),
    .INIT_58(256'h000000108200130000000032b680b2020000001cf502065e0000000b203206a2),
    .INIT_59(256'h00000022b613656400000011f011c32000000013a0011301000000139002071c),
    .INIT_5A(256'h000000118012254200000032b70206600000001cf302066400000001f0020684),
    .INIT_5B(256'h00000022b692004700000011f012003e000000138002065e000000139002068e),
    .INIT_5C(256'h0000000b0132005000000003a03325780000002f9111d0020000002f8100b002),
    .INIT_5D(256'h0000002fa122005900000004a0032578000000140061d003000000140060b002),
    .INIT_5E(256'h0000001d000200470000000b0132003e0000002500022587000000370002085b),
    .INIT_5F(256'h0000001d03020050000000030f0325840000000b0391d00200000032b810b002),
    .INIT_60(256'h00000020b9e2005900000022b843258400000020b971d00300000032b830b002),
    .INIT_61(256'h000000096080100000000009508206c60000002f50301060000000095082085b),
    .INIT_62(256'h000000096080100000000009508207000000002f6052d0030000002f5042f032),
    .INIT_63(256'h0000000960801d00000000095082200a0000002f631207130000002f530206d2),
    .INIT_64(256'h000000096082fe11000000095082fd100000002f63801f000000002f53701e00),
    .INIT_65(256'h000000015ef2fd13000000250002fd010000002f60601d000000002f53c2ff12),
    .INIT_66(256'h0000002d60a0b00f0000002d50920ba5000000011002fd1e0000000160701d01),
    .INIT_67(256'h0000000160b03007000000015c30b00f00000025000325ba0000002d10b1d0ff),
    .INIT_68(256'h0000002d10b325aa0000002d60a1d0000000002d5090b001000000011002f00f),
    .INIT_69(256'h0000000b810325b200000020b7a1d00200000037001325ae000000250001d001),
    .INIT_6A(256'h0000002f935207cd0000002f834208e80000000ba12325b60000000b9111d003),
    .INIT_6B(256'h0000000b330207d40000000bd37208eb00000001200221720000002fa362093c),
    .INIT_6C(256'h0000001ba00207de0000001a940208ee00000018830221720000000b4312093c),
    .INIT_6D(256'h0000002f935207ea0000002f834208f100000011201221720000003abbc2093c),
    .INIT_6E(256'h00000022bb10d00400000032be80900e0000001c2d0221720000002fa362093c),
    .INIT_6F(256'h0000002f20f2b04e0000000ba362f0330000000b935090160000000b834325c3),
    .INIT_70(256'h0000001d4010b00400000009408325e4000000013001d00e000000012000300f),
    .INIT_71(256'h0000001ba000be110000001b9000bd10000000188400b20600000032c7a0b105),
    .INIT_72(256'h0000002f8341ee10000000133001cd000000001120103f030000003abcf0bf12),
    .INIT_73(256'h0000000b83413e0000000022bc211d010000002fa36325d50000002f9351ef20),
    .INIT_74(256'h0000002f20d2ff120000002f30e2fe110000000ba362fd100000000b93513f00),
    .INIT_75(256'h0000000b60e191010000000b50d0b1020000000b40c0b0010000002f80c22598),
    .INIT_76(256'h000000146082f00100000014608110010000000b30e325e40000000b70f1c010),
    .INIT_77(256'h0000002f70e01f000000001470001e000000001430801d00000000147002f013),
    .INIT_78(256'h0000001400622598000000140062ff12000000140062fe110000000b0132fd10),
    .INIT_79(256'h000000250000100000000037000207af0000002f00f20037000000140062079f),
    .INIT_7A(256'h00000032c1e207130000001d400206d2000000034f0010000000000b4392d003),
    .INIT_7B(256'h0000001b900365ed000000188400d080000000012000900d0000000b43c2200a),
    .INIT_7C(256'h0000002f834365f1000000112010d0400000003abf90900d0000001ba0025000),
    .INIT_7D(256'h00000032c1e205f10000001d2022df070000002fa36205f10000002f93525000),
    .INIT_7E(256'h0000000ba36205f10000000b9352dd070000000b834205f100000022bee2de07),
    .INIT_7F(256'h00000018840205f1000000194022db070000000b43c205f10000002f20f2dc07),
    .INITP_00(256'hb8be8abe9dbe0d3a19b48c89829fb109a48da60623b30824141c991ab6038f12),
    .INITP_01(256'h1dbb071d9e8335982410bb84a8bb9ea39e8b1792bb101a9d2f81a79a360c3b02),
    .INITP_02(256'ha53f240226bf0ab30e9882929ea738063e83bb01bf982216bd2210bb01b99824),
    .INITP_03(256'h87bca4a323ba05ad8ea181ba06ba0604a22c158416289d859e92159e1a8b0310),
    .INITP_04(256'h271f21a711b99f0285b531b5abb83090af8590823b353729ac3e152f09009489),
    .INITP_05(256'hba901634b503021a98a00926119636a8bf26a61c0224021eba3bb38a3f9436ac),
    .INITP_06(256'ha793180fa4353a3903982106b58c1ba6348e8326a534118fac882abf339d1ba4),
    .INITP_07(256'h1b13228b279513869925b7b8b6b3839ca93c0f298b0e258606328e9430b7afa0),
    .INITP_08(256'hadba94b62b180d891d319b0509303683bd061d08b52bb8279f8b010333293a2e),
    .INITP_09(256'hb830041d8a10a3a6a038140a3d87320bb7950232ae033a20b5123b278a090802),
    .INITP_0A(256'h290682ac259828a9b18d22989eb4ac07229302b9b21204bf150da599043f35b7),
    .INITP_0B(256'h9b97a32713aaa82436b406142f1321890002123fb839bc3f028c22b203b28395),
    .INITP_0C(256'h3b30bfb11c0f8db9b6a5a7a01c1b32b81010ae3a030d252b0384b4933a812fbc),
    .INITP_0D(256'h8833aa0f898c952d369ab68f1d822212b013072d3c973ea7872ba924230a1e94),
    .INITP_0E(256'h17a219388a992399a1a496839930ac2d19a9bfb186a7282282859f9622ae2105),
    .INITP_0F(256'h140e129eb3b08c37ba29b63318aa249d009986063cb73a84303b349c01838837),
