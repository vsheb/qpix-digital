    .INIT_00(256'h00000020a512f01e00000020a330100000000020a272b80f0000000b92f2b40f),
    .INIT_01(256'h00000014b002070200000014a0e207690000000ba252f03200000001b0001001),
    .INIT_02(256'h00000014a00206dc00000014b002247a00000014a00206de0000000ba26206e2),
    .INIT_03(256'h0000000b21d2b80f00000014b002b40f00000014a002b20f00000014b0020896),
    .INIT_04(256'h00000014b00224bb00000014a00207690000002f21d2f032000000062b001002),
    .INIT_05(256'h00000014b00206b600000014a000bc0b00000014b00206de00000014a0020716),
    .INIT_06(256'h00000014b00206b600000014a000bc0900000014b00206b600000014a000bc0a),
    .INIT_07(256'h00000014a00206b600000014b000bc0700000014a00206b60000000ba270bc08),
    .INIT_08(256'h0000000b21c3242800000014b000d00800000014a000900200000014b00206dc),
    .INIT_09(256'h00000001a0022008000000250002074d0000002fb1c0101000000006b2020896),
    .INIT_0A(256'h0000000d8ff2200800000014a002077b0000000d1ff2074d00000001b0001000),
    .INIT_0B(256'h0000000daff0bd0a00000014a000bc090000000d9ff0bb0800000014a000ba07),
    .INIT_0C(256'h00000000200030f000000025000000e00000002fb2501f0000000014b000be0b),
    .INIT_0D(256'h00000014a043243900000014a000d0800000000d1ff3243900000001a001d0c0),
    .INIT_0E(256'h00000014a042f01400000014a040301f00000014a04000a000000014a0422475),
    .INIT_0F(256'h000000022a0000b000000014a04206a200000014a04206a200000014a04206a2),
    .INIT_10(256'h000000250002f0150000002f2263e475000000062b01d07b00000020a440307f),
    .INIT_11(256'h00000014b00000f000000014a062f01300000000b900300300000000a80000e0),
    .INIT_12(256'h00000014b002fd1100000014a062fc1000000014b00206a200000014a0603003),
    .INIT_13(256'h00000014b002f01300000014a063645f00000014b000df0800000014a062fe12),
    .INIT_14(256'h00000001a001cab0000000003800bb02000000002100ba130000002500003f01),
    .INIT_15(256'h0000000d2ff2fe0e000000033012fd0d000000032aa2fc0c00000001b0036475),
    .INIT_16(256'h0000000daff03f0300000014a0014f000000000d3ff14e0600000014a002ff0f),
    .INIT_17(256'h00000001a000ba130000000038022472000000002103247500000014b081df01),
    .INIT_18(256'h00000014a0003e010000000d2ff36475000000033021cab0000000032cc0bb02),
    .INIT_19(256'h00000014b080b0040000000daff2fe1200000014a002fd110000000d3ff2fc10),
    .INIT_1A(256'h000000032f01ad1000000001a0018c00000000003800b206000000002100b105),
    .INIT_1B(256'h0000000d3ff0b40f00000014a0020b5f0000000d2ff3e475000000033041ae20),
    .INIT_1C(256'h0000002fb272068700000014b08208fa0000000daff2f40f00000014a0003401),
    .INIT_1D(256'h0000000100c2074d000000008400100000000000950208a500000025000208fe),
    .INIT_1E(256'h000000131000d040000000148080900f0000001490e22008000000011002077b),
    .INIT_1F(256'h00000036a830d0800000001d1003618b00000036a790d020000000190013618b),
    .INIT_20(256'h0000000d50836182000000250000d080000000018ff0900e000000019ff36186),
    .INIT_21(256'h000000018ff3617c000000019ff0d020000000011023617f00000036a890d040),
    .INIT_22(256'h000000001500d0040000003ea950900e0000001d10336179000000250000d010),
    .INIT_23(256'h0000001410e2b04e000000118012f00b000000018ff0901b0000000004032494),
    .INIT_24(256'h000000011042247a0000000190f324a30000003ea8e1d0e000000014008030f0),
    .INIT_25(256'h0000001982809006000000008403647a000000009500d020000000250000900d),
    .INIT_26(256'h000000019ff3647a000000011021d0530000003ea9e324a30000001b9041d049),
    .INIT_27(256'h0000000381f20702000000001802078400000025000206dc000000018ff20720),
    .INIT_28(256'h000000149002070c000000141062247a00000014900206de00000014106206e2),
    .INIT_29(256'h0000001d90f208a5000000011022012d000000149002089600000014106206dc),
    .INIT_2A(256'h0000000110401000000000390002d0030000001d80c2f03200000036aab01000),
    .INIT_2B(256'h0000000b20c2089600000020b4622008000000370012077b000000250002074d),
    .INIT_2C(256'h00000014206207410000000ba0f010600000000b40e208a50000000b30d2012d),
    .INIT_2D(256'h000000142080100000000014a002d003000000144002f0320000001430001000),
    .INIT_2E(256'h0000001450e01d000000000340322008000000005402077b0000000327f2074d),
    .INIT_2F(256'h000000007a02fe11000000036032fd10000000006a001f000000001450e01e00),
    .INIT_30(256'h00000001d0020b5f000000037032fd1e0000001470e01d010000001470e2ff12),
    .INIT_31(256'h00000032aea0b00f0000001d602324cd000000008201d0ff00000001e000b00f),
    .INIT_32(256'h00000001a002091100000001900208fa00000032b112f00f0000001d60303001),
    .INIT_33(256'h00000032ad7324d60000001ce400d00400000036ad00900e0000001cd30221ad),
    .INIT_34(256'h00000013a00030f0000000139002b04e000000108f02f00b00000009f080901b),
    .INIT_35(256'h00000001d000b10500000022acc0b00400000013e00324e800000011d011d0e0),
    .INIT_36(256'h00000032ae10bf120000001cd500be110000000bf310bd100000000be300b206),
    .INIT_37(256'h00000011d011ef2000000013a001ee10000000129f01cd00000000108e003f01),
    .INIT_38(256'h00000003a0113f000000002f91113e000000002f81011d0100000022ada324e8),
    .INIT_39(256'h0000002fa12224c100000004a002ff12000000140062fe110000000b0022fd10),
    .INIT_3A(256'h0000000be31010000000000bd30208a5000000250002012d0000003700020896),
    .INIT_3B(256'h00000001f002077b00000001a002074d00000001900010000000000b2372d103),
    .INIT_3C(256'h000000129e03654b000000108d01d00100000032af70b01e0000001cf2022008),
    .INIT_3D(256'h00000001f0020a7500000022af00b51700000011f010b41600000013a0001200),
    .INIT_3E(256'h000000108200b41800000032b00042100000001cf502f9170000000b23c2f816),
    .INIT_3F(256'h00000022af92f91900000011f012f81800000013a0020a75000000139000b519),
    .INIT_40(256'h0000001180220a7500000032b080b51b0000001cf300b41a00000001f0004210),
    .INIT_41(256'h00000022b010b41c00000011f0104210000000138002f91b000000139002f81a),
    .INIT_42(256'h0000000b0022f91d00000003a012f81c0000002f91120a750000002f8100b51d),
    .INIT_43(256'h00000037000012020000002fa123251c00000004a000d2020000001400604210),
    .INIT_44(256'h0000000b237208110000000be31208040000000bd3020819000000250002f21e),
    .INIT_45(256'h00000001f001d00200000001a00324af000000019001d001000000018000b032),
    .INIT_46(256'h000000129e02258c000000108d00502000000032b1f2073b0000001cf20324cd),
    .INIT_47(256'h0000000bf390b01600000022b1820c1500000011f012f21e00000013a0001204),
    .INIT_48(256'h00000001f001d0ff00000032b2c2f1150000001df002f01400000003ff00b117),
    .INIT_49(256'h000000108200b11900000032b2c0b0180000001df02346870000000b23c1f1ff),
    .INIT_4A(256'h00000022b251f1ff00000011f011d0ff00000013a002f115000000139002f014),
    .INIT_4B(256'h00000032b352f0140000001cf500b11b0000000b2380b01a00000001f0034687),
    .INIT_4C(256'h00000011f013468700000013a001f1ff000000139001d0ff000000108202f115),
    .INIT_4D(256'h00000032b3d2f1150000001cf302f01400000001f000b11d00000022b2e0b01c),
    .INIT_4E(256'h00000011f010b0320000001380034687000000139001f1ff000000118011d0ff),
    .INIT_4F(256'h00000003a01208190000002f911208fe0000002f8103653f00000022b361d000),
    .INIT_50(256'h0000002fa120b03200000004a002081100000014006208400000000b00220804),
    .INIT_51(256'h00000009508324cd00000020b581d00200000025000324af000000370001d001),
    .INIT_52(256'h000000095081d0080000002f6052258c0000002f504030df000000096082073b),
    .INIT_53(256'h00000009508207000000002f6312071e0000002f530207000000000960836558),
    .INIT_54(256'h000000095081d0010000002f6380b0320000002f537207e900000009608206dc),
    .INIT_55(256'h000000250002258c0000002f606050200000002f53c2073b00000009608324af),
    .INIT_56(256'h0000002d5092072400000001100206fc0000000160736565000000015f01d010),
    .INIT_57(256'h000000370010b03200000025000207e90000002d10b206dc0000002d60a2072a),
    .INIT_58(256'h0000000ba12050200000000b9112073b0000000b810324af00000020b461d001),
    .INIT_59(256'h00000001200206fc0000002fa36365720000002f9351d0200000002f8342258c),
    .INIT_5A(256'h00000018830207e90000000b431206dc0000000b3302072a0000000bd3720724),
    .INIT_5B(256'h000000112012073b0000003ab76324af0000001ba001d0010000001a9400b032),
    .INIT_5C(256'h0000001c2d03657f0000002fa361d0400000002f9352258c0000002f834030df),
    .INIT_5D(256'h0000000b935206dc0000000b8342072a00000022b6b2072400000032ba8206fc),
    .INIT_5E(256'h00000001300324af000000012001d0010000002f20f0b0320000000ba36207e9),
    .INIT_5F(256'h000000188401d08000000032c0e2258c0000001d401030df000000094082073b),
    .INIT_60(256'h00000011201207140000003ab89207180000001ba002071e0000001b90036017),
    .INIT_61(256'h0000002fa361d0010000002f9350b0320000002f834207e900000013300206dc),
    .INIT_62(256'h0000000ba362258c0000000b935030df0000000b8342073b00000022b7c324af),
    .INIT_63(256'h0000000b40c220080000002f80c2074d0000002f20d010080000002f30e20741),
    .INIT_64(256'h00000014408090020000001450836604000000144061d0040000000b50d0b01e),
    .INIT_65(256'h00000014608206760000000b60e206500000000b50d325ef0000002f40c0d004),
    .INIT_66(256'h0000000b70f1ff320000000b60e1dedb0000002f50d0bf05000000145080be04),
    .INIT_67(256'h0000000377f011bb0000001470001ed00000001460801f0900000014608325a2),
    .INIT_68(256'h0000001400601e400000000b00201f0a00000001700225a60000002f70e0120b),
    .INIT_69(256'h0000002500009d0700000037000206280000002f70f0120c000000047000112b),
    .INIT_6A(256'h00000032bdf1ce100000001d4002dd08000000034f02de090000000b4392df0a),
    .INIT_6B(256'h0000001b900225b300000018840365b0000000012001cf200000000b43c365b0),
    .INIT_6C(256'h0000002f8340b01600000011201225a60000003abb913f000000001ba0011e01),
    .INIT_6D(256'h00000032bdf1d0ff0000001d2022f1150000002fa362f0140000002f9350b117),
    .INIT_6E(256'h0000000ba36012000000000b935206300000000b834325bf00000022bae1f1ff),
    .INIT_6F(256'h000000188400b018000000194022f2200000000b43c142000000002f20f0d0ff),
    .INIT_70(256'h0000000b8341d0ff0000003ec0e2f1150000001ba002f0140000001b9000b119),
    .INIT_71(256'h00000000380012000000000b20f206300000000ba36325cb0000000b9351f1ff),
    .INIT_72(256'h000000143060b01a000000148082f2210000001490e14200000000033010d0ff),
    .INIT_73(256'h000000148061d0ff0000002f30c2f115000000143082f014000000148080b11b),
    .INIT_74(256'h00000014908012000000002f80d2063000000014808325d7000000149081f1ff),
    .INIT_75(256'h0000002f20e0b01c0000001420e2f2220000001420614200000000142000d0ff),
    .INIT_76(256'h000000043002f115000000140062f0140000000b00201200000000013010b11d),
    .INIT_77(256'h0000000b4382063000000025000325e4000000370001f1ff0000002f30f1d0ff),
    .INIT_78(256'h0000001ba002f2230000001b90014200000000188400d0ff0000000120001200),
    .INIT_79(256'h0000002f9350b0200000002f8342081100000011201208590000003abea2080c),
    .INIT_7A(256'h0000000b935040100000000b8340b12200000022be1040100000002fa360b121),
    .INIT_7B(256'h000000194022073b0000000b438325f20000002f20f040100000000ba360b123),
    .INIT_7C(256'h0000003ec0e030bf0000001ba002073b0000001b900225f40000001884005040),
    .INIT_7D(256'h0000000b20f0b01f0000000ba362f03b0000000b9350b00e0000000b83420741),
    .INIT_7E(256'h0000002f30c2b20f00000014308208a500000014808366000000000b30019001),
    .INIT_7F(256'h0000002f80d226250000001480801002000000149082b80f000000148062b40f),
    .INITP_00(256'h9a299aa8b90eb908b98b3f91a61e901191288a2399a21ca1bd04af17913c3934),
    .INITP_01(256'h3e89898984931a1a869f9fa7a1af17a6a10e228b83121794a6b0853f0e3702ba),
    .INITP_02(256'ha1a32a253e9f300d01141882a2a6bebd3b0b2a0cad87b600a79f1a2db98d0a1d),
    .INITP_03(256'h38aababa9f391e9634153f2419be3b8d3d00131ea338bca6ac2f8ea1120694aa),
    .INITP_04(256'h29903b92239e951d0684a32719bf1e1ab7a60c3f89172a3881b99bb93d3d80a4),
    .INITP_05(256'h9202b31c1f28b5992982b69732b41f2b0028a9b00a88b9b70f0d87bf1da79bb8),
    .INITP_06(256'h253b008e2e39349a1b96143e23ad999bbd3b9a8424a21a0da48d3f13872538bc),
    .INITP_07(256'h051a23ba079d110d269b03ba9496abb0313730128b81b0a1a82d88b31d268c8a),
    .INITP_08(256'hb923863c119c09aba3b9249391998fb6b8bf33163e99a4052c8101acb48dbd30),
    .INITP_09(256'h9c279826801ab936823531bc0a3ea784910202bb24943039060a889925061399),
    .INITP_0A(256'ha9302e1c1e97bbafa9aa3f0d90afa8080dacbc9014ac32888eaf3e27b5a7083e),
    .INITP_0B(256'h8f3d382cbc8596333e8d90bd9aaaa993ab9f8a9fb402300e10ad2d902ebd012d),
    .INITP_0C(256'h9cac950d0aa4311b832a22113818a3a102958a2eaaaf871822b009baa6149a84),
    .INITP_0D(256'h1c8b8c943db2869a15263c3285b18a1b040d030b1dbab81db63a9f9f8cb30605),
    .INITP_0E(256'h0939b9a1b89d222802aa2d368688a702253000281da91182b99437bf9823941f),
    .INITP_0F(256'h172e0f28ac9dbeb01b34370dbc158f0b810d99b4ba083e34bc97b2391907169f),
