    .INIT_00(256'h0250003240501f010207ec1d0032ff0000bc0c0b00201f0000bd0d202b228000),
    .INIT_01(256'h0207be2243601001001101010022003300108020766280000207ef202bb2df02),
    .INIT_02(256'h0207ec2200a2df020207dc2057601f0000110001082320770010002f01f20560),
    .INIT_03(256'h0207a0324272202a0207f21d0082202a025000324272202a0207031d00228000),
    .INIT_04(256'h001004364192202a0207be1d0202202a001101324272202a0010801d0102202a),
    .INIT_05(256'h02070f010022202a0207ec205542202a0207dc050402202a0011002054b2202a),
    .INIT_06(256'h0010802054b2202a0207a6364202202a0207f51d0402202a025000224362202a),
    .INIT_07(256'h0011002243628000001008010022df020207be2055401f01001101030bf2202a),
    .INIT_08(256'h025000030bf1d0040207202054b320770207ec3602a1d0010207dc1d0802054e),
    .INIT_09(256'h0011012027120551001080224363239b0207b0010021d0080207f820554322c4),
    .INIT_0A(256'h0207dc32431205540011001d0020106000100c0b002322c40207be2027a1d004),
    .INIT_0B(256'h00900e32431205220250001d0032051a0207350b002205600207ec202830109f),
    .INIT_0C(256'h00900e05040200370250002054b22bfc03682f20766204ec00d0082028c20532),
    .INIT_0D(256'h00900f2058e090020250002056025000032833010002006300d002205542004a),
    .INIT_0E(256'h009010364390d0010250000d0800b0000328370900d3204600d0022200a0d080),
    .INIT_0F(256'h0090113643d0121f0250000d040011ff03283b0900d010ff00d0022500036046),
    .INIT_10(256'h000950013003e0400250000150a1b20003283f014401b10000d0022500019001),
    .INIT_11(256'h01490e142000d0400011000d0100900100100c0b0142f0000008400b21501001),
    .INIT_12(256'h036847143002b00c019001142002b0000131000d008250000148081430032046),
    .INIT_13(256'h0018ff3a4522d0100019ff19001010ff036851011012bfff01d100030072bf7e),
    .INIT_14(256'h001102123502d001036857102400300f00d5082244e09001025000141062d011),
    .INIT_15(256'h01d103020100900602500009008360590018ff2d2090d0200019ff2d30a0900d),
    .INIT_16(256'h0018ff14b060900d0000400bb130900600015001a000900603e8642500022054),
    .INIT_17(256'h03e85c09e1e2205b01400809d1d0900701410e09c1c3606001180114b060d080),
    .INIT_18(256'h02500013d002053000110410cb02500000190b10ba00900701180809f1f09007),
    .INIT_19(256'h01b90501b002053401981801a04204f000084013f002052400095013e0020514),
    .INIT_1A(256'h0018ff204392050c0019ff09c072052e001102204392053203e86d2048320522),
    .INIT_1B(256'h01410620439204f000381f09e07204f6000180204392053602500009d07204f0),
    .INIT_1C(256'h0141060b4100101901490001b012500001410601a73204ec01490009f07204f4),
    .INIT_1D(256'h000a9010c402021900008003601250000011020b6123e0740149000b51119001),
    .INIT_1E(256'h01400619a010d00101400613f000900d01400612e602020701400612d5020221),
    .INIT_1F(256'h01da5d01a7401080014a0025000206b10140063e477206aa014a001bb003207a),
    .INIT_20(256'h01d8142043d1dc9303688525000207e901d90b20483207be03d00001b0101101),
    .INIT_21(256'h01d8082043d207d50250002de07010000011042043d0110003a8872df073607d),
    .INIT_22(256'h0095082043d1d11202089e2dc070311e0250002043d001e003a8852dd072088a),
    .INIT_23(256'h02f504250001d1160096082da07320a00095082043d1d11402f5032db0732092),
    .INIT_24(256'h02f5300b2152f2390096080130001220009508015002202a02f6050146c320ac),
    .INIT_25(256'h02f5371430014008009608142001410a0095080d010001e002f6310b014000d0),
    .INIT_26(256'h02f53c030071d04800960814300320b8009508142001d05802f6380d008030f8),
    .INIT_27(256'h001607141062202a0015ef3a4a1320bb025000190011d08802f60601101320b8),
    .INIT_28(256'h02d10b2d30a001e002d60a12350000d002d509102402f2390011002249d01220),
    .INIT_29(256'h00b1172d30a1d04800b01606010030f800130009008140080250002d2091410a),
    .INIT_2A(256'h02f22014a062202a02f11725000320be02f0162d0081d0880208c22d209320bb),
    .INIT_2B(256'h0208c214e00001e000b11914d00000d000b01814c002f23900130114b0001230),
    .INIT_2C(256'h00130214e081d08802f22114f0e030f802f119250001400802f01814f001410a),
    .INIT_2D(256'h02f01a14a082202a0208c214b08320bb00b11b14c081d0c800b01a14d08320b8),
    .INIT_2E(256'h00b01c190e90100300130339000220c002f222110b92f00202f11b2500001002),
    .INIT_2F(256'h02f11d110072f00202f01c3e4c3010040208c219011220c000b11d390002f002),
    .INIT_30(256'h01d0ff1100a01000001200250002f201025000190f60120302f2233900020203),
    .INIT_31(256'h014006204d720213014006204cd2f02403100000c000100101f1ff250002f03a),
    .INIT_32(256'h0140062054020235014100204d72022c014006204cd20247014006205402023e),
    .INIT_33(256'h01400e141000101001400e14c060110001400e01100207e90141002500020266),
    .INIT_34(256'h022bfc141000110002500014c060101000b224141002026601003014c06207d5),
    .INIT_35(256'h022bfc1d10a207d5022bfc2500001010022bfc1410001100022bfc14c0620250),
    .INIT_36(256'h022bfc25000206aa022bfc1113020760022bfc11107206aa022bfc3a4da20792),
    .INIT_37(256'h022bfc204b9207e9022bfc09006207be022bfc2054301101022bfc01a0001080),
    .INIT_38(256'h022bfc19101207a0022bfc204ab207d5022bfc0110401004022bfc3900001100),
    .INIT_39(256'h022bfc204d7207a0022bfc0010020235022bfc04a00207a0022bfc364e22022c),
    .INIT_3A(256'h022bfc25000206aa022bfc364dd20247022bfc19201207a0022bfc205402023e),
    .INIT_3B(256'h022bfc22540207e9022bfc0112020266022bfc22540206aa022bfc0110d20760),
    .INIT_3C(256'h022bfc22540010c0022bfc0113e207d5022bfc2254001014022bfc0115f01100),
    .INIT_3D(256'h022bfc2254001014022bfc01133207a0022bfc22540207be022bfc0113101101),
    .INIT_3E(256'h022bfc2254001014022bfc0113101100022bfc2254020250022bfc0113001100),
    .INIT_3F(256'h022bfc2254032159022bfc011331d002022bfc225400b002022bfc01132207d5),
    .INIT_40(256'h022bfc22540206aa022bfc0113520760022bfc22540206aa022bfc0113420792),
    .INIT_41(256'h022bfc2254001101022bfc0113701080022bfc22540206aa022bfc0113620760),
    .INIT_42(256'h022bfc2254001008022bfc0113901100022bfc22540207e9022bfc01138207be),
    .INIT_43(256'h022bfc22540207a6022bfc011422022c022bfc22540207a6022bfc01141207d5),
    .INIT_44(256'h022bfc22540207a6022bfc011442023e022bfc22540207a6022bfc0114320235),
    .INIT_45(256'h022bfc22540206aa022bfc0114620760022bfc22540206aa022bfc0114520247),
    .INIT_46(256'h022bfc22540207e9022bfc0114820266022bfc22540206aa022bfc0114720760),
    .INIT_47(256'h022bfc22540010c0022bfc0114a207d5022bfc2254001018022bfc0114901100),
    .INIT_48(256'h022bfc2254001018022bfc0114c207a6022bfc22540207be022bfc0114b01101),
    .INIT_49(256'h022bfc2254001018022bfc0114e01100022bfc2254020250022bfc0114d01100),
    .INIT_4A(256'h022bfc2254032159022bfc011501d003022bfc225400b002022bfc0114f207d5),
    .INIT_4B(256'h022bfc22540206aa022bfc0115220760022bfc22540206aa022bfc0115120792),
    .INIT_4C(256'h022bfc22540206aa022bfc0115420760022bfc22540206aa022bfc0115320760),
    .INIT_4D(256'h022bfc22540207e9022bfc01156207be022bfc2254001101022bfc0115501080),
    .INIT_4E(256'h022bfc22540207b0022bfc01158207d5022bfc225400100c022bfc0115701100),
    .INIT_4F(256'h022bfc22540207b0022bfc0115a20235022bfc22540207b0022bfc011592022c),
    .INIT_50(256'h022bfc0900d206aa022bfc2500020247022bfc2d106207b0022bfc205472023e),
    .INIT_51(256'h022bfc0900d206aa022bfc2500020760022bfc36543206aa022bfc0d02020760),
    .INIT_52(256'h022bfc09000207e9022bfc2500020266022bfc36547206aa022bfc0d01020760),
    .INIT_53(256'h022bfc0309f010c0022bfc09000207d5022bfc250000101c022bfc0306001100),
    .INIT_54(256'h022bfc250000101c022bfc03007207b0022bfc09013207be022bfc2500001101),
    .INIT_55(256'h022bfc041000101c022bfc2054e01100022bfc0316020250022bfc0010001100),
    .INIT_56(256'h022bfc204ee207a0022bfc20510206b4022bfc20516206b7022bfc2d100207d5),
    .INIT_57(256'h022bfc250000b002022bfc204ec206b4022bfc204c5207a0022bfc2054b206b7),
    .INIT_58(256'h022bfc04100206b7022bfc2054b207a6022bfc0319f3216d022bfc001001d002),
    .INIT_59(256'h022bfc204ee1d003022bfc205100b002022bfc20530206b4022bfc2d100207a6),
    .INIT_5A(256'h022bfc2054e207b0022bfc3258a206b7022bfc1d001207b0022bfc0b0323216d),
    .INIT_5B(256'h022bfc205300b002022bfc25000202a9022bfc204ec202a0022bfc204c5206b4),
    .INIT_5C(256'h022bfc204c50b002022bfc01002202b2022bfc204ee32177022bfc205101d002),
    .INIT_5D(256'h022bfc0319f20766022bfc00100202bb022bfc2500032177022bfc204ec1d003),
    .INIT_5E(256'h022bfc2500001002022bfc2d1002d00f022bfc0410001002022bfc2054b2b02e),
    .INIT_5F(256'h022bfc2d10320833022bfc0b1322d011022bfc2057601002022bfc010002d010),
    .INIT_60(256'h022bfc0b0322d00f022bfc204ee01002022bfc2051020837022bfc205302b02e),
    .INIT_61(256'h022bfc204c52083b022bfc0104032190022bfc3258a1d002022bfc1d0010b002),
    .INIT_62(256'h022bfc204c51d003022bfc010200b002022bfc250002d010022bfc204ec01002),
    .INIT_63(256'h022bfc1d0002d011022bfc2054e01002022bfc250002083f022bfc204ec32190),
    .INIT_64(256'h022bfc204ee01002022bfc204f220837022bfc205282b02e022bfc3259520833),
    .INIT_65(256'h022bfc20530321a1022bfc225921d002022bfc2051c0b002022bfc250002d00f),
    .INIT_66(256'h022bfc204c60b002022bfc00c302d010022bfc204ee01002022bfc205262083b),
    .INIT_67(256'h022bfc2052e01002022bfc205592083f022bfc20565321a1022bfc204ec1d003),
    .INIT_68(256'h022bfc204c62020d022bfc0bc3a20203022bfc204ee20792022bfc2051c2d011),
    .INIT_69(256'h022bfc2051601100022bfc2052401010022bfc2500020266022bfc204ec206aa),
    .INIT_6A(256'h022bfc0bc06207d5022bfc204f801010022bfc204f801100022bfc204ee2025b),
    .INIT_6B(256'h022bfc0bc0401100022bfc204c601014022bfc0bc0520266022bfc204c6207a0),
    .INIT_6C(256'h022bfc20532207d5022bfc205fc01014022bfc204ec01100022bfc204c62025b),
    .INIT_6D(256'h022bfc0d504207a6022bfc09502321ca022bfc204ee1d002022bfc2050e0b002),
    .INIT_6E(256'h022bfc09c1c2025b022bfc225d201100022bfc2060e01018022bfc3a5bb20266),
    .INIT_6F(256'h022bfc0bb130b002022bfc09f1f207d5022bfc09e1e01018022bfc09d1d01100),
    .INIT_70(256'h022bfc13d0020266022bfc10cb0207b0022bfc14b06321ca022bfc14b061d003),
    .INIT_71(256'h022bfc2fe3601100022bfc2ff3b2025b022bfc13f0001100022bfc13e000101c),
    .INIT_72(256'h022bfc204c62b04e022bfc0bc3b20203022bfc2fc34207d5022bfc2fd350101c),
    .INIT_73(256'h022bfc204c6321f1022bfc0bc351d001022bfc204c60300f022bfc0bc3609001),
    .INIT_74(256'h022bfc2051020766022bfc204ec321e2022bfc204c60d002022bfc0bc3409002),
    .INIT_75(256'h022bfc3a5da2b04f022bfc0d5042b80f022bfc204ee2b40f022bfc2050e2b20f),
    .INIT_76(256'h022bfc0bd352d010022bfc0bc34010e0022bfc225f02b10f022bfc2060e2b08f),
    .INIT_77(256'h022bfc01b0020560022bfc01a0401002022bfc0bf3b2d010022bfc0be360101c),
    .INIT_78(256'h022bfc204392027a022bfc09f0720271022bfc204392200a022bfc204832058e),
    .INIT_79(256'h022bfc2043920283022bfc09d07321ec022bfc204391d002022bfc09e070b002),
    .INIT_7A(256'h022bfc204c62028c022bfc00cd0321ec022bfc204c61d003022bfc09c070b002),
    .INIT_7B(256'h022bfc204c62058e022bfc00cf020560022bfc204c601000022bfc00ce020766),
    .INIT_7C(256'h022bfc204ee2b40f022bfc205222b20f022bfc2051020766022bfc204ec2200a),
    .INIT_7D(256'h022bfc14c002b10f022bfc0d5042b08f022bfc01c002b04f022bfc204f82b80f),
    .INIT_7E(256'h022bfc250002d010022bfc204ec0101c022bfc204c62d010022bfc11c01010e0),
    .INIT_7F(256'h022bfc2b80c20512022bfc204ee2057c022bfc205302f032022bfc2053201001),
    .INITP_00(256'h2929f08396c4cfec5bc66717bc692790f15dc3feddc68811438db877c7478813),
    .INITP_01(256'h325ed5240355dd9509c2d79f8d43ce323d57c4f8448b1bd885bf785568ceda73),
    .INITP_02(256'hd71f102ab8aa90e99dd7ab2200459a6f1003ef30d9b0a79582320807b3eccf38),
    .INITP_03(256'h28b825372da6008f1ab380ba35822481a73a9b6b022620e6032436925527ab9c),
    .INITP_04(256'hbe8575c1d4a91f4a629d83c54b809472dab5adf2aedad4d30ce7b1c3b4dd1d46),
    .INITP_05(256'h6e6a690920a243d9656a09adb278fbcfed8ca7a742d4ec7f9396a1616a4fda1c),
    .INITP_06(256'h70d559747f7b6f6f75f6715271da3e2e8ba8270c172e80161c0957a007bb7e43),
    .INITP_07(256'hf54b7dc1f1cf77d5f1d6fc4c7940f16bfecffeca7f78ca5a5bf3f9794df7c3da),
    .INITP_08(256'h797c7072feecfe6dfe77fe7e72e8727472637260f952fe4770c9fe57fed6fecd),
    .INITP_09(256'hf86df8e1f8797ff6fee370ecfe72feeffef5fe75f5f77d7a70ef776e70f5fc6a),
    .INITP_0A(256'hfcc45ec15de465f4df41c6f377494df169d2776150f6e1efcb77fd6ecbfff7c7),
    .INITP_0B(256'h66ddd5e5fae75255c67bfad852e0577bf5f6445c4adbce6c43eafbfa5cc643ec),
    .INITP_0C(256'h775fc7d8d3c057f9feea6bee57da6a5fcec96f4140e6e0cc47d3424b73577e69),
    .INITP_0D(256'hc5c8fd78c454e468efc5c06e6ffb44d8ea5f74dffe42c65ae37df6495971dbf4),
    .INITP_0E(256'hdd617e51c06bc6f058e44bf562cc54f65a68c46bce6be152516cf0d6d05071e8),
    .INITP_0F(256'hf8dcf56ee041cfc547f9644c4b6b62dd5f5a50c956c2c14d536cc0e953c946f8),
